library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_buzzer is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant buzzer_lut : array_1d := (
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    1    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    2    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    3    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    4    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    5    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    6    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    7    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    8    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    9    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    10    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    11    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    12    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    13    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    14    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    15    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    16    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    17    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    18    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    19    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )    ,
   (    20    )   
);

end package LUT_buzzer;
