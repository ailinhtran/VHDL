library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_ledr is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant ledr_LUT : array_1d := (
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	511	)	,
    (	510	)	,
    (	510	)	,
    (	510	)	,
    (	510	)	,
    (	510	)	,
    (	510	)	,
    (	510	)	,
    (	509	)	,
    (	509	)	,
    (	509	)	,
    (	509	)	,
    (	509	)	,
    (	509	)	,
    (	509	)	,
    (	509	)	,
    (	508	)	,
    (	508	)	,
    (	508	)	,
    (	508	)	,
    (	508	)	,
    (	508	)	,
    (	508	)	,
    (	507	)	,
    (	507	)	,
    (	507	)	,
    (	507	)	,
    (	507	)	,
    (	507	)	,
    (	507	)	,
    (	506	)	,
    (	506	)	,
    (	506	)	,
    (	506	)	,
    (	506	)	,
    (	506	)	,
    (	506	)	,
    (	505	)	,
    (	505	)	,
    (	505	)	,
    (	505	)	,
    (	505	)	,
    (	505	)	,
    (	505	)	,
    (	505	)	,
    (	504	)	,
    (	504	)	,
    (	504	)	,
    (	504	)	,
    (	504	)	,
    (	504	)	,
    (	504	)	,
    (	503	)	,
    (	503	)	,
    (	503	)	,
    (	503	)	,
    (	503	)	,
    (	503	)	,
    (	503	)	,
    (	502	)	,
    (	502	)	,
    (	502	)	,
    (	502	)	,
    (	502	)	,
    (	502	)	,
    (	502	)	,
    (	501	)	,
    (	501	)	,
    (	501	)	,
    (	501	)	,
    (	501	)	,
    (	501	)	,
    (	501	)	,
    (	501	)	,
    (	500	)	,
    (	500	)	,
    (	500	)	,
    (	500	)	,
    (	500	)	,
    (	500	)	,
    (	500	)	,
    (	499	)	,
    (	499	)	,
    (	499	)	,
    (	499	)	,
    (	499	)	,
    (	499	)	,
    (	499	)	,
    (	498	)	,
    (	498	)	,
    (	498	)	,
    (	498	)	,
    (	498	)	,
    (	498	)	,
    (	498	)	,
    (	497	)	,
    (	497	)	,
    (	497	)	,
    (	497	)	,
    (	497	)	,
    (	497	)	,
    (	497	)	,
    (	497	)	,
    (	496	)	,
    (	496	)	,
    (	496	)	,
    (	496	)	,
    (	496	)	,
    (	496	)	,
    (	496	)	,
    (	495	)	,
    (	495	)	,
    (	495	)	,
    (	495	)	,
    (	495	)	,
    (	495	)	,
    (	495	)	,
    (	494	)	,
    (	494	)	,
    (	494	)	,
    (	494	)	,
    (	494	)	,
    (	494	)	,
    (	494	)	,
    (	493	)	,
    (	493	)	,
    (	493	)	,
    (	493	)	,
    (	493	)	,
    (	493	)	,
    (	493	)	,
    (	492	)	,
    (	492	)	,
    (	492	)	,
    (	492	)	,
    (	492	)	,
    (	492	)	,
    (	492	)	,
    (	492	)	,
    (	491	)	,
    (	491	)	,
    (	491	)	,
    (	491	)	,
    (	491	)	,
    (	491	)	,
    (	491	)	,
    (	490	)	,
    (	490	)	,
    (	490	)	,
    (	490	)	,
    (	490	)	,
    (	490	)	,
    (	490	)	,
    (	489	)	,
    (	489	)	,
    (	489	)	,
    (	489	)	,
    (	489	)	,
    (	489	)	,
    (	489	)	,
    (	488	)	,
    (	488	)	,
    (	488	)	,
    (	488	)	,
    (	488	)	,
    (	488	)	,
    (	488	)	,
    (	488	)	,
    (	487	)	,
    (	487	)	,
    (	487	)	,
    (	487	)	,
    (	487	)	,
    (	487	)	,
    (	487	)	,
    (	486	)	,
    (	486	)	,
    (	486	)	,
    (	486	)	,
    (	486	)	,
    (	486	)	,
    (	486	)	,
    (	485	)	,
    (	485	)	,
    (	485	)	,
    (	485	)	,
    (	485	)	,
    (	485	)	,
    (	485	)	,
    (	484	)	,
    (	484	)	,
    (	484	)	,
    (	484	)	,
    (	484	)	,
    (	484	)	,
    (	484	)	,
    (	484	)	,
    (	483	)	,
    (	483	)	,
    (	483	)	,
    (	483	)	,
    (	483	)	,
    (	483	)	,
    (	483	)	,
    (	482	)	,
    (	482	)	,
    (	482	)	,
    (	482	)	,
    (	482	)	,
    (	482	)	,
    (	482	)	,
    (	481	)	,
    (	481	)	,
    (	481	)	,
    (	481	)	,
    (	481	)	,
    (	481	)	,
    (	481	)	,
    (	480	)	,
    (	480	)	,
    (	480	)	,
    (	480	)	,
    (	480	)	,
    (	480	)	,
    (	480	)	,
    (	480	)	,
    (	479	)	,
    (	479	)	,
    (	479	)	,
    (	479	)	,
    (	479	)	,
    (	479	)	,
    (	479	)	,
    (	478	)	,
    (	478	)	,
    (	478	)	,
    (	478	)	,
    (	478	)	,
    (	478	)	,
    (	478	)	,
    (	477	)	,
    (	477	)	,
    (	477	)	,
    (	477	)	,
    (	477	)	,
    (	477	)	,
    (	477	)	,
    (	476	)	,
    (	476	)	,
    (	476	)	,
    (	476	)	,
    (	476	)	,
    (	476	)	,
    (	476	)	,
    (	476	)	,
    (	475	)	,
    (	475	)	,
    (	475	)	,
    (	475	)	,
    (	475	)	,
    (	475	)	,
    (	475	)	,
    (	474	)	,
    (	474	)	,
    (	474	)	,
    (	474	)	,
    (	474	)	,
    (	474	)	,
    (	474	)	,
    (	473	)	,
    (	473	)	,
    (	473	)	,
    (	473	)	,
    (	473	)	,
    (	473	)	,
    (	473	)	,
    (	472	)	,
    (	472	)	,
    (	472	)	,
    (	472	)	,
    (	472	)	,
    (	472	)	,
    (	472	)	,
    (	472	)	,
    (	471	)	,
    (	471	)	,
    (	471	)	,
    (	471	)	,
    (	471	)	,
    (	471	)	,
    (	471	)	,
    (	470	)	,
    (	470	)	,
    (	470	)	,
    (	470	)	,
    (	470	)	,
    (	470	)	,
    (	470	)	,
    (	469	)	,
    (	469	)	,
    (	469	)	,
    (	469	)	,
    (	469	)	,
    (	469	)	,
    (	469	)	,
    (	468	)	,
    (	468	)	,
    (	468	)	,
    (	468	)	,
    (	468	)	,
    (	468	)	,
    (	468	)	,
    (	468	)	,
    (	467	)	,
    (	467	)	,
    (	467	)	,
    (	467	)	,
    (	467	)	,
    (	467	)	,
    (	467	)	,
    (	466	)	,
    (	466	)	,
    (	466	)	,
    (	466	)	,
    (	466	)	,
    (	466	)	,
    (	466	)	,
    (	465	)	,
    (	465	)	,
    (	465	)	,
    (	465	)	,
    (	465	)	,
    (	465	)	,
    (	465	)	,
    (	464	)	,
    (	464	)	,
    (	464	)	,
    (	464	)	,
    (	464	)	,
    (	464	)	,
    (	464	)	,
    (	464	)	,
    (	463	)	,
    (	463	)	,
    (	463	)	,
    (	463	)	,
    (	463	)	,
    (	463	)	,
    (	463	)	,
    (	462	)	,
    (	462	)	,
    (	462	)	,
    (	462	)	,
    (	462	)	,
    (	462	)	,
    (	462	)	,
    (	461	)	,
    (	461	)	,
    (	461	)	,
    (	461	)	,
    (	461	)	,
    (	461	)	,
    (	461	)	,
    (	460	)	,
    (	460	)	,
    (	460	)	,
    (	460	)	,
    (	460	)	,
    (	460	)	,
    (	460	)	,
    (	459	)	,
    (	459	)	,
    (	459	)	,
    (	459	)	,
    (	459	)	,
    (	459	)	,
    (	459	)	,
    (	459	)	,
    (	458	)	,
    (	458	)	,
    (	458	)	,
    (	458	)	,
    (	458	)	,
    (	458	)	,
    (	458	)	,
    (	457	)	,
    (	457	)	,
    (	457	)	,
    (	457	)	,
    (	457	)	,
    (	457	)	,
    (	457	)	,
    (	456	)	,
    (	456	)	,
    (	456	)	,
    (	456	)	,
    (	456	)	,
    (	456	)	,
    (	456	)	,
    (	455	)	,
    (	455	)	,
    (	455	)	,
    (	455	)	,
    (	455	)	,
    (	455	)	,
    (	455	)	,
    (	455	)	,
    (	454	)	,
    (	454	)	,
    (	454	)	,
    (	454	)	,
    (	454	)	,
    (	454	)	,
    (	454	)	,
    (	453	)	,
    (	453	)	,
    (	453	)	,
    (	453	)	,
    (	453	)	,
    (	453	)	,
    (	453	)	,
    (	452	)	,
    (	452	)	,
    (	452	)	,
    (	452	)	,
    (	452	)	,
    (	452	)	,
    (	452	)	,
    (	451	)	,
    (	451	)	,
    (	451	)	,
    (	451	)	,
    (	451	)	,
    (	451	)	,
    (	451	)	,
    (	451	)	,
    (	450	)	,
    (	450	)	,
    (	450	)	,
    (	450	)	,
    (	450	)	,
    (	450	)	,
    (	450	)	,
    (	449	)	,
    (	449	)	,
    (	449	)	,
    (	449	)	,
    (	449	)	,
    (	449	)	,
    (	449	)	,
    (	448	)	,
    (	448	)	,
    (	448	)	,
    (	448	)	,
    (	448	)	,
    (	448	)	,
    (	448	)	,
    (	447	)	,
    (	447	)	,
    (	447	)	,
    (	447	)	,
    (	447	)	,
    (	447	)	,
    (	447	)	,
    (	447	)	,
    (	446	)	,
    (	446	)	,
    (	446	)	,
    (	446	)	,
    (	446	)	,
    (	446	)	,
    (	446	)	,
    (	445	)	,
    (	445	)	,
    (	445	)	,
    (	445	)	,
    (	445	)	,
    (	445	)	,
    (	445	)	,
    (	444	)	,
    (	444	)	,
    (	444	)	,
    (	444	)	,
    (	444	)	,
    (	444	)	,
    (	444	)	,
    (	443	)	,
    (	443	)	,
    (	443	)	,
    (	443	)	,
    (	443	)	,
    (	443	)	,
    (	443	)	,
    (	443	)	,
    (	442	)	,
    (	442	)	,
    (	442	)	,
    (	442	)	,
    (	442	)	,
    (	442	)	,
    (	442	)	,
    (	441	)	,
    (	441	)	,
    (	441	)	,
    (	441	)	,
    (	441	)	,
    (	441	)	,
    (	441	)	,
    (	440	)	,
    (	440	)	,
    (	440	)	,
    (	440	)	,
    (	440	)	,
    (	440	)	,
    (	440	)	,
    (	439	)	,
    (	439	)	,
    (	439	)	,
    (	439	)	,
    (	439	)	,
    (	439	)	,
    (	439	)	,
    (	439	)	,
    (	438	)	,
    (	438	)	,
    (	438	)	,
    (	438	)	,
    (	438	)	,
    (	438	)	,
    (	438	)	,
    (	437	)	,
    (	437	)	,
    (	437	)	,
    (	437	)	,
    (	437	)	,
    (	437	)	,
    (	437	)	,
    (	436	)	,
    (	436	)	,
    (	436	)	,
    (	436	)	,
    (	436	)	,
    (	436	)	,
    (	436	)	,
    (	435	)	,
    (	435	)	,
    (	435	)	,
    (	435	)	,
    (	435	)	,
    (	435	)	,
    (	435	)	,
    (	435	)	,
    (	434	)	,
    (	434	)	,
    (	434	)	,
    (	434	)	,
    (	434	)	,
    (	434	)	,
    (	434	)	,
    (	433	)	,
    (	433	)	,
    (	433	)	,
    (	433	)	,
    (	433	)	,
    (	433	)	,
    (	433	)	,
    (	432	)	,
    (	432	)	,
    (	432	)	,
    (	432	)	,
    (	432	)	,
    (	432	)	,
    (	432	)	,
    (	431	)	,
    (	431	)	,
    (	431	)	,
    (	431	)	,
    (	431	)	,
    (	431	)	,
    (	431	)	,
    (	431	)	,
    (	430	)	,
    (	430	)	,
    (	430	)	,
    (	430	)	,
    (	430	)	,
    (	430	)	,
    (	430	)	,
    (	429	)	,
    (	429	)	,
    (	429	)	,
    (	429	)	,
    (	429	)	,
    (	429	)	,
    (	429	)	,
    (	428	)	,
    (	428	)	,
    (	428	)	,
    (	428	)	,
    (	428	)	,
    (	428	)	,
    (	428	)	,
    (	427	)	,
    (	427	)	,
    (	427	)	,
    (	427	)	,
    (	427	)	,
    (	427	)	,
    (	427	)	,
    (	427	)	,
    (	426	)	,
    (	426	)	,
    (	426	)	,
    (	426	)	,
    (	426	)	,
    (	426	)	,
    (	426	)	,
    (	425	)	,
    (	425	)	,
    (	425	)	,
    (	425	)	,
    (	425	)	,
    (	425	)	,
    (	425	)	,
    (	424	)	,
    (	424	)	,
    (	424	)	,
    (	424	)	,
    (	424	)	,
    (	424	)	,
    (	424	)	,
    (	423	)	,
    (	423	)	,
    (	423	)	,
    (	423	)	,
    (	423	)	,
    (	423	)	,
    (	423	)	,
    (	422	)	,
    (	422	)	,
    (	422	)	,
    (	422	)	,
    (	422	)	,
    (	422	)	,
    (	422	)	,
    (	422	)	,
    (	421	)	,
    (	421	)	,
    (	421	)	,
    (	421	)	,
    (	421	)	,
    (	421	)	,
    (	421	)	,
    (	420	)	,
    (	420	)	,
    (	420	)	,
    (	420	)	,
    (	420	)	,
    (	420	)	,
    (	420	)	,
    (	419	)	,
    (	419	)	,
    (	419	)	,
    (	419	)	,
    (	419	)	,
    (	419	)	,
    (	419	)	,
    (	418	)	,
    (	418	)	,
    (	418	)	,
    (	418	)	,
    (	418	)	,
    (	418	)	,
    (	418	)	,
    (	418	)	,
    (	417	)	,
    (	417	)	,
    (	417	)	,
    (	417	)	,
    (	417	)	,
    (	417	)	,
    (	417	)	,
    (	416	)	,
    (	416	)	,
    (	416	)	,
    (	416	)	,
    (	416	)	,
    (	416	)	,
    (	416	)	,
    (	415	)	,
    (	415	)	,
    (	415	)	,
    (	415	)	,
    (	415	)	,
    (	415	)	,
    (	415	)	,
    (	414	)	,
    (	414	)	,
    (	414	)	,
    (	414	)	,
    (	414	)	,
    (	414	)	,
    (	414	)	,
    (	414	)	,
    (	413	)	,
    (	413	)	,
    (	413	)	,
    (	413	)	,
    (	413	)	,
    (	413	)	,
    (	413	)	,
    (	412	)	,
    (	412	)	,
    (	412	)	,
    (	412	)	,
    (	412	)	,
    (	412	)	,
    (	412	)	,
    (	411	)	,
    (	411	)	,
    (	411	)	,
    (	411	)	,
    (	411	)	,
    (	411	)	,
    (	411	)	,
    (	410	)	,
    (	410	)	,
    (	410	)	,
    (	410	)	,
    (	410	)	,
    (	410	)	,
    (	410	)	,
    (	410	)	,
    (	409	)	,
    (	409	)	,
    (	409	)	,
    (	409	)	,
    (	409	)	,
    (	409	)	,
    (	409	)	,
    (	408	)	,
    (	408	)	,
    (	408	)	,
    (	408	)	,
    (	408	)	,
    (	408	)	,
    (	408	)	,
    (	407	)	,
    (	407	)	,
    (	407	)	,
    (	407	)	,
    (	407	)	,
    (	407	)	,
    (	407	)	,
    (	406	)	,
    (	406	)	,
    (	406	)	,
    (	406	)	,
    (	406	)	,
    (	406	)	,
    (	406	)	,
    (	406	)	,
    (	405	)	,
    (	405	)	,
    (	405	)	,
    (	405	)	,
    (	405	)	,
    (	405	)	,
    (	405	)	,
    (	404	)	,
    (	404	)	,
    (	404	)	,
    (	404	)	,
    (	404	)	,
    (	404	)	,
    (	404	)	,
    (	403	)	,
    (	403	)	,
    (	403	)	,
    (	403	)	,
    (	403	)	,
    (	403	)	,
    (	403	)	,
    (	402	)	,
    (	402	)	,
    (	402	)	,
    (	402	)	,
    (	402	)	,
    (	402	)	,
    (	402	)	,
    (	402	)	,
    (	401	)	,
    (	401	)	,
    (	401	)	,
    (	401	)	,
    (	401	)	,
    (	401	)	,
    (	401	)	,
    (	400	)	,
    (	400	)	,
    (	400	)	,
    (	400	)	,
    (	400	)	,
    (	400	)	,
    (	400	)	,
    (	399	)	,
    (	399	)	,
    (	399	)	,
    (	399	)	,
    (	399	)	,
    (	399	)	,
    (	399	)	,
    (	398	)	,
    (	398	)	,
    (	398	)	,
    (	398	)	,
    (	398	)	,
    (	398	)	,
    (	398	)	,
    (	398	)	,
    (	397	)	,
    (	397	)	,
    (	397	)	,
    (	397	)	,
    (	397	)	,
    (	397	)	,
    (	397	)	,
    (	396	)	,
    (	396	)	,
    (	396	)	,
    (	396	)	,
    (	396	)	,
    (	396	)	,
    (	396	)	,
    (	395	)	,
    (	395	)	,
    (	395	)	,
    (	395	)	,
    (	395	)	,
    (	395	)	,
    (	395	)	,
    (	394	)	,
    (	394	)	,
    (	394	)	,
    (	394	)	,
    (	394	)	,
    (	394	)	,
    (	394	)	,
    (	394	)	,
    (	393	)	,
    (	393	)	,
    (	393	)	,
    (	393	)	,
    (	393	)	,
    (	393	)	,
    (	393	)	,
    (	392	)	,
    (	392	)	,
    (	392	)	,
    (	392	)	,
    (	392	)	,
    (	392	)	,
    (	392	)	,
    (	391	)	,
    (	391	)	,
    (	391	)	,
    (	391	)	,
    (	391	)	,
    (	391	)	,
    (	391	)	,
    (	390	)	,
    (	390	)	,
    (	390	)	,
    (	390	)	,
    (	390	)	,
    (	390	)	,
    (	390	)	,
    (	389	)	,
    (	389	)	,
    (	389	)	,
    (	389	)	,
    (	389	)	,
    (	389	)	,
    (	389	)	,
    (	389	)	,
    (	388	)	,
    (	388	)	,
    (	388	)	,
    (	388	)	,
    (	388	)	,
    (	388	)	,
    (	388	)	,
    (	387	)	,
    (	387	)	,
    (	387	)	,
    (	387	)	,
    (	387	)	,
    (	387	)	,
    (	387	)	,
    (	386	)	,
    (	386	)	,
    (	386	)	,
    (	386	)	,
    (	386	)	,
    (	386	)	,
    (	386	)	,
    (	385	)	,
    (	385	)	,
    (	385	)	,
    (	385	)	,
    (	385	)	,
    (	385	)	,
    (	385	)	,
    (	385	)	,
    (	384	)	,
    (	384	)	,
    (	384	)	,
    (	384	)	,
    (	384	)	,
    (	384	)	,
    (	384	)	,
    (	383	)	,
    (	383	)	,
    (	383	)	,
    (	383	)	,
    (	383	)	,
    (	383	)	,
    (	383	)	,
    (	382	)	,
    (	382	)	,
    (	382	)	,
    (	382	)	,
    (	382	)	,
    (	382	)	,
    (	382	)	,
    (	381	)	,
    (	381	)	,
    (	381	)	,
    (	381	)	,
    (	381	)	,
    (	381	)	,
    (	381	)	,
    (	381	)	,
    (	380	)	,
    (	380	)	,
    (	380	)	,
    (	380	)	,
    (	380	)	,
    (	380	)	,
    (	380	)	,
    (	379	)	,
    (	379	)	,
    (	379	)	,
    (	379	)	,
    (	379	)	,
    (	379	)	,
    (	379	)	,
    (	378	)	,
    (	378	)	,
    (	378	)	,
    (	378	)	,
    (	378	)	,
    (	378	)	,
    (	378	)	,
    (	377	)	,
    (	377	)	,
    (	377	)	,
    (	377	)	,
    (	377	)	,
    (	377	)	,
    (	377	)	,
    (	377	)	,
    (	376	)	,
    (	376	)	,
    (	376	)	,
    (	376	)	,
    (	376	)	,
    (	376	)	,
    (	376	)	,
    (	375	)	,
    (	375	)	,
    (	375	)	,
    (	375	)	,
    (	375	)	,
    (	375	)	,
    (	375	)	,
    (	374	)	,
    (	374	)	,
    (	374	)	,
    (	374	)	,
    (	374	)	,
    (	374	)	,
    (	374	)	,
    (	373	)	,
    (	373	)	,
    (	373	)	,
    (	373	)	,
    (	373	)	,
    (	373	)	,
    (	373	)	,
    (	373	)	,
    (	372	)	,
    (	372	)	,
    (	372	)	,
    (	372	)	,
    (	372	)	,
    (	372	)	,
    (	372	)	,
    (	371	)	,
    (	371	)	,
    (	371	)	,
    (	371	)	,
    (	371	)	,
    (	371	)	,
    (	371	)	,
    (	370	)	,
    (	370	)	,
    (	370	)	,
    (	370	)	,
    (	370	)	,
    (	370	)	,
    (	370	)	,
    (	369	)	,
    (	369	)	,
    (	369	)	,
    (	369	)	,
    (	369	)	,
    (	369	)	,
    (	369	)	,
    (	369	)	,
    (	368	)	,
    (	368	)	,
    (	368	)	,
    (	368	)	,
    (	368	)	,
    (	368	)	,
    (	368	)	,
    (	367	)	,
    (	367	)	,
    (	367	)	,
    (	367	)	,
    (	367	)	,
    (	367	)	,
    (	367	)	,
    (	366	)	,
    (	366	)	,
    (	366	)	,
    (	366	)	,
    (	366	)	,
    (	366	)	,
    (	366	)	,
    (	365	)	,
    (	365	)	,
    (	365	)	,
    (	365	)	,
    (	365	)	,
    (	365	)	,
    (	365	)	,
    (	365	)	,
    (	364	)	,
    (	364	)	,
    (	364	)	,
    (	364	)	,
    (	364	)	,
    (	364	)	,
    (	364	)	,
    (	363	)	,
    (	363	)	,
    (	363	)	,
    (	363	)	,
    (	363	)	,
    (	363	)	,
    (	363	)	,
    (	362	)	,
    (	362	)	,
    (	362	)	,
    (	362	)	,
    (	362	)	,
    (	362	)	,
    (	362	)	,
    (	361	)	,
    (	361	)	,
    (	361	)	,
    (	361	)	,
    (	361	)	,
    (	361	)	,
    (	361	)	,
    (	361	)	,
    (	360	)	,
    (	360	)	,
    (	360	)	,
    (	360	)	,
    (	360	)	,
    (	360	)	,
    (	360	)	,
    (	359	)	,
    (	359	)	,
    (	359	)	,
    (	359	)	,
    (	359	)	,
    (	359	)	,
    (	359	)	,
    (	358	)	,
    (	358	)	,
    (	358	)	,
    (	358	)	,
    (	358	)	,
    (	358	)	,
    (	358	)	,
    (	357	)	,
    (	357	)	,
    (	357	)	,
    (	357	)	,
    (	357	)	,
    (	357	)	,
    (	357	)	,
    (	356	)	,
    (	356	)	,
    (	356	)	,
    (	356	)	,
    (	356	)	,
    (	356	)	,
    (	356	)	,
    (	356	)	,
    (	355	)	,
    (	355	)	,
    (	355	)	,
    (	355	)	,
    (	355	)	,
    (	355	)	,
    (	355	)	,
    (	354	)	,
    (	354	)	,
    (	354	)	,
    (	354	)	,
    (	354	)	,
    (	354	)	,
    (	354	)	,
    (	353	)	,
    (	353	)	,
    (	353	)	,
    (	353	)	,
    (	353	)	,
    (	353	)	,
    (	353	)	,
    (	352	)	,
    (	352	)	,
    (	352	)	,
    (	352	)	,
    (	352	)	,
    (	352	)	,
    (	352	)	,
    (	352	)	,
    (	351	)	,
    (	351	)	,
    (	351	)	,
    (	351	)	,
    (	351	)	,
    (	351	)	,
    (	351	)	,
    (	350	)	,
    (	350	)	,
    (	350	)	,
    (	350	)	,
    (	350	)	,
    (	350	)	,
    (	350	)	,
    (	349	)	,
    (	349	)	,
    (	349	)	,
    (	349	)	,
    (	349	)	,
    (	349	)	,
    (	349	)	,
    (	348	)	,
    (	348	)	,
    (	348	)	,
    (	348	)	,
    (	348	)	,
    (	348	)	,
    (	348	)	,
    (	348	)	,
    (	347	)	,
    (	347	)	,
    (	347	)	,
    (	347	)	,
    (	347	)	,
    (	347	)	,
    (	347	)	,
    (	346	)	,
    (	346	)	,
    (	346	)	,
    (	346	)	,
    (	346	)	,
    (	346	)	,
    (	346	)	,
    (	345	)	,
    (	345	)	,
    (	345	)	,
    (	345	)	,
    (	345	)	,
    (	345	)	,
    (	345	)	,
    (	344	)	,
    (	344	)	,
    (	344	)	,
    (	344	)	,
    (	344	)	,
    (	344	)	,
    (	344	)	,
    (	344	)	,
    (	343	)	,
    (	343	)	,
    (	343	)	,
    (	343	)	,
    (	343	)	,
    (	343	)	,
    (	343	)	,
    (	342	)	,
    (	342	)	,
    (	342	)	,
    (	342	)	,
    (	342	)	,
    (	342	)	,
    (	342	)	,
    (	341	)	,
    (	341	)	,
    (	341	)	,
    (	341	)	,
    (	341	)	,
    (	341	)	,
    (	341	)	,
    (	340	)	,
    (	340	)	,
    (	340	)	,
    (	340	)	,
    (	340	)	,
    (	340	)	,
    (	340	)	,
    (	340	)	,
    (	339	)	,
    (	339	)	,
    (	339	)	,
    (	339	)	,
    (	339	)	,
    (	339	)	,
    (	339	)	,
    (	338	)	,
    (	338	)	,
    (	338	)	,
    (	338	)	,
    (	338	)	,
    (	338	)	,
    (	338	)	,
    (	337	)	,
    (	337	)	,
    (	337	)	,
    (	337	)	,
    (	337	)	,
    (	337	)	,
    (	337	)	,
    (	336	)	,
    (	336	)	,
    (	336	)	,
    (	336	)	,
    (	336	)	,
    (	336	)	,
    (	336	)	,
    (	336	)	,
    (	335	)	,
    (	335	)	,
    (	335	)	,
    (	335	)	,
    (	335	)	,
    (	335	)	,
    (	335	)	,
    (	334	)	,
    (	334	)	,
    (	334	)	,
    (	334	)	,
    (	334	)	,
    (	334	)	,
    (	334	)	,
    (	333	)	,
    (	333	)	,
    (	333	)	,
    (	333	)	,
    (	333	)	,
    (	333	)	,
    (	333	)	,
    (	332	)	,
    (	332	)	,
    (	332	)	,
    (	332	)	,
    (	332	)	,
    (	332	)	,
    (	332	)	,
    (	332	)	,
    (	331	)	,
    (	331	)	,
    (	331	)	,
    (	331	)	,
    (	331	)	,
    (	331	)	,
    (	331	)	,
    (	330	)	,
    (	330	)	,
    (	330	)	,
    (	330	)	,
    (	330	)	,
    (	330	)	,
    (	330	)	,
    (	329	)	,
    (	329	)	,
    (	329	)	,
    (	329	)	,
    (	329	)	,
    (	329	)	,
    (	329	)	,
    (	328	)	,
    (	328	)	,
    (	328	)	,
    (	328	)	,
    (	328	)	,
    (	328	)	,
    (	328	)	,
    (	328	)	,
    (	327	)	,
    (	327	)	,
    (	327	)	,
    (	327	)	,
    (	327	)	,
    (	327	)	,
    (	327	)	,
    (	326	)	,
    (	326	)	,
    (	326	)	,
    (	326	)	,
    (	326	)	,
    (	326	)	,
    (	326	)	,
    (	325	)	,
    (	325	)	,
    (	325	)	,
    (	325	)	,
    (	325	)	,
    (	325	)	,
    (	325	)	,
    (	324	)	,
    (	324	)	,
    (	324	)	,
    (	324	)	,
    (	324	)	,
    (	324	)	,
    (	324	)	,
    (	323	)	,
    (	323	)	,
    (	323	)	,
    (	323	)	,
    (	323	)	,
    (	323	)	,
    (	323	)	,
    (	323	)	,
    (	322	)	,
    (	322	)	,
    (	322	)	,
    (	322	)	,
    (	322	)	,
    (	322	)	,
    (	322	)	,
    (	321	)	,
    (	321	)	,
    (	321	)	,
    (	321	)	,
    (	321	)	,
    (	321	)	,
    (	321	)	,
    (	320	)	,
    (	320	)	,
    (	320	)	,
    (	320	)	,
    (	320	)	,
    (	320	)	,
    (	320	)	,
    (	319	)	,
    (	319	)	,
    (	319	)	,
    (	319	)	,
    (	319	)	,
    (	319	)	,
    (	319	)	,
    (	319	)	,
    (	318	)	,
    (	318	)	,
    (	318	)	,
    (	318	)	,
    (	318	)	,
    (	318	)	,
    (	318	)	,
    (	317	)	,
    (	317	)	,
    (	317	)	,
    (	317	)	,
    (	317	)	,
    (	317	)	,
    (	317	)	,
    (	316	)	,
    (	316	)	,
    (	316	)	,
    (	316	)	,
    (	316	)	,
    (	316	)	,
    (	316	)	,
    (	315	)	,
    (	315	)	,
    (	315	)	,
    (	315	)	,
    (	315	)	,
    (	315	)	,
    (	315	)	,
    (	315	)	,
    (	314	)	,
    (	314	)	,
    (	314	)	,
    (	314	)	,
    (	314	)	,
    (	314	)	,
    (	314	)	,
    (	313	)	,
    (	313	)	,
    (	313	)	,
    (	313	)	,
    (	313	)	,
    (	313	)	,
    (	313	)	,
    (	312	)	,
    (	312	)	,
    (	312	)	,
    (	312	)	,
    (	312	)	,
    (	312	)	,
    (	312	)	,
    (	311	)	,
    (	311	)	,
    (	311	)	,
    (	311	)	,
    (	311	)	,
    (	311	)	,
    (	311	)	,
    (	311	)	,
    (	310	)	,
    (	310	)	,
    (	310	)	,
    (	310	)	,
    (	310	)	,
    (	310	)	,
    (	310	)	,
    (	309	)	,
    (	309	)	,
    (	309	)	,
    (	309	)	,
    (	309	)	,
    (	309	)	,
    (	309	)	,
    (	308	)	,
    (	308	)	,
    (	308	)	,
    (	308	)	,
    (	308	)	,
    (	308	)	,
    (	308	)	,
    (	307	)	,
    (	307	)	,
    (	307	)	,
    (	307	)	,
    (	307	)	,
    (	307	)	,
    (	307	)	,
    (	307	)	,
    (	306	)	,
    (	306	)	,
    (	306	)	,
    (	306	)	,
    (	306	)	,
    (	306	)	,
    (	306	)	,
    (	305	)	,
    (	305	)	,
    (	305	)	,
    (	305	)	,
    (	305	)	,
    (	305	)	,
    (	305	)	,
    (	304	)	,
    (	304	)	,
    (	304	)	,
    (	304	)	,
    (	304	)	,
    (	304	)	,
    (	304	)	,
    (	303	)	,
    (	303	)	,
    (	303	)	,
    (	303	)	,
    (	303	)	,
    (	303	)	,
    (	303	)	,
    (	303	)	,
    (	302	)	,
    (	302	)	,
    (	302	)	,
    (	302	)	,
    (	302	)	,
    (	302	)	,
    (	302	)	,
    (	301	)	,
    (	301	)	,
    (	301	)	,
    (	301	)	,
    (	301	)	,
    (	301	)	,
    (	301	)	,
    (	300	)	,
    (	300	)	,
    (	300	)	,
    (	300	)	,
    (	300	)	,
    (	300	)	,
    (	300	)	,
    (	299	)	,
    (	299	)	,
    (	299	)	,
    (	299	)	,
    (	299	)	,
    (	299	)	,
    (	299	)	,
    (	299	)	,
    (	298	)	,
    (	298	)	,
    (	298	)	,
    (	298	)	,
    (	298	)	,
    (	298	)	,
    (	298	)	,
    (	297	)	,
    (	297	)	,
    (	297	)	,
    (	297	)	,
    (	297	)	,
    (	297	)	,
    (	297	)	,
    (	296	)	,
    (	296	)	,
    (	296	)	,
    (	296	)	,
    (	296	)	,
    (	296	)	,
    (	296	)	,
    (	295	)	,
    (	295	)	,
    (	295	)	,
    (	295	)	,
    (	295	)	,
    (	295	)	,
    (	295	)	,
    (	295	)	,
    (	294	)	,
    (	294	)	,
    (	294	)	,
    (	294	)	,
    (	294	)	,
    (	294	)	,
    (	294	)	,
    (	293	)	,
    (	293	)	,
    (	293	)	,
    (	293	)	,
    (	293	)	,
    (	293	)	,
    (	293	)	,
    (	292	)	,
    (	292	)	,
    (	292	)	,
    (	292	)	,
    (	292	)	,
    (	292	)	,
    (	292	)	,
    (	291	)	,
    (	291	)	,
    (	291	)	,
    (	291	)	,
    (	291	)	,
    (	291	)	,
    (	291	)	,
    (	291	)	,
    (	290	)	,
    (	290	)	,
    (	290	)	,
    (	290	)	,
    (	290	)	,
    (	290	)	,
    (	290	)	,
    (	289	)	,
    (	289	)	,
    (	289	)	,
    (	289	)	,
    (	289	)	,
    (	289	)	,
    (	289	)	,
    (	288	)	,
    (	288	)	,
    (	288	)	,
    (	288	)	,
    (	288	)	,
    (	288	)	,
    (	288	)	,
    (	287	)	,
    (	287	)	,
    (	287	)	,
    (	287	)	,
    (	287	)	,
    (	287	)	,
    (	287	)	,
    (	286	)	,
    (	286	)	,
    (	286	)	,
    (	286	)	,
    (	286	)	,
    (	286	)	,
    (	286	)	,
    (	286	)	,
    (	285	)	,
    (	285	)	,
    (	285	)	,
    (	285	)	,
    (	285	)	,
    (	285	)	,
    (	285	)	,
    (	284	)	,
    (	284	)	,
    (	284	)	,
    (	284	)	,
    (	284	)	,
    (	284	)	,
    (	284	)	,
    (	283	)	,
    (	283	)	,
    (	283	)	,
    (	283	)	,
    (	283	)	,
    (	283	)	,
    (	283	)	,
    (	282	)	,
    (	282	)	,
    (	282	)	,
    (	282	)	,
    (	282	)	,
    (	282	)	,
    (	282	)	,
    (	282	)	,
    (	281	)	,
    (	281	)	,
    (	281	)	,
    (	281	)	,
    (	281	)	,
    (	281	)	,
    (	281	)	,
    (	280	)	,
    (	280	)	,
    (	280	)	,
    (	280	)	,
    (	280	)	,
    (	280	)	,
    (	280	)	,
    (	279	)	,
    (	279	)	,
    (	279	)	,
    (	279	)	,
    (	279	)	,
    (	279	)	,
    (	279	)	,
    (	278	)	,
    (	278	)	,
    (	278	)	,
    (	278	)	,
    (	278	)	,
    (	278	)	,
    (	278	)	,
    (	278	)	,
    (	277	)	,
    (	277	)	,
    (	277	)	,
    (	277	)	,
    (	277	)	,
    (	277	)	,
    (	277	)	,
    (	276	)	,
    (	276	)	,
    (	276	)	,
    (	276	)	,
    (	276	)	,
    (	276	)	,
    (	276	)	,
    (	275	)	,
    (	275	)	,
    (	275	)	,
    (	275	)	,
    (	275	)	,
    (	275	)	,
    (	275	)	,
    (	274	)	,
    (	274	)	,
    (	274	)	,
    (	274	)	,
    (	274	)	,
    (	274	)	,
    (	274	)	,
    (	274	)	,
    (	273	)	,
    (	273	)	,
    (	273	)	,
    (	273	)	,
    (	273	)	,
    (	273	)	,
    (	273	)	,
    (	272	)	,
    (	272	)	,
    (	272	)	,
    (	272	)	,
    (	272	)	,
    (	272	)	,
    (	272	)	,
    (	271	)	,
    (	271	)	,
    (	271	)	,
    (	271	)	,
    (	271	)	,
    (	271	)	,
    (	271	)	,
    (	270	)	,
    (	270	)	,
    (	270	)	,
    (	270	)	,
    (	270	)	,
    (	270	)	,
    (	270	)	,
    (	270	)	,
    (	269	)	,
    (	269	)	,
    (	269	)	,
    (	269	)	,
    (	269	)	,
    (	269	)	,
    (	269	)	,
    (	268	)	,
    (	268	)	,
    (	268	)	,
    (	268	)	,
    (	268	)	,
    (	268	)	,
    (	268	)	,
    (	267	)	,
    (	267	)	,
    (	267	)	,
    (	267	)	,
    (	267	)	,
    (	267	)	,
    (	267	)	,
    (	266	)	,
    (	266	)	,
    (	266	)	,
    (	266	)	,
    (	266	)	,
    (	266	)	,
    (	266	)	,
    (	266	)	,
    (	265	)	,
    (	265	)	,
    (	265	)	,
    (	265	)	,
    (	265	)	,
    (	265	)	,
    (	265	)	,
    (	264	)	,
    (	264	)	,
    (	264	)	,
    (	264	)	,
    (	264	)	,
    (	264	)	,
    (	264	)	,
    (	263	)	,
    (	263	)	,
    (	263	)	,
    (	263	)	,
    (	263	)	,
    (	263	)	,
    (	263	)	,
    (	262	)	,
    (	262	)	,
    (	262	)	,
    (	262	)	,
    (	262	)	,
    (	262	)	,
    (	262	)	,
    (	262	)	,
    (	261	)	,
    (	261	)	,
    (	261	)	,
    (	261	)	,
    (	261	)	,
    (	261	)	,
    (	261	)	,
    (	260	)	,
    (	260	)	,
    (	260	)	,
    (	260	)	,
    (	260	)	,
    (	260	)	,
    (	260	)	,
    (	259	)	,
    (	259	)	,
    (	259	)	,
    (	259	)	,
    (	259	)	,
    (	259	)	,
    (	259	)	,
    (	258	)	,
    (	258	)	,
    (	258	)	,
    (	258	)	,
    (	258	)	,
    (	258	)	,
    (	258	)	,
    (	258	)	,
    (	257	)	,
    (	257	)	,
    (	257	)	,
    (	257	)	,
    (	257	)	,
    (	257	)	,
    (	257	)	,
    (	256	)	,
    (	256	)	,
    (	256	)	,
    (	256	)	,
    (	256	)	,
    (	256	)	,
    (	256	)	,
    (	255	)	,
    (	255	)	,
    (	255	)	,
    (	255	)	,
    (	255	)	,
    (	255	)	,
    (	255	)	,
    (	254	)	,
    (	254	)	,
    (	254	)	,
    (	254	)	,
    (	254	)	,
    (	254	)	,
    (	254	)	,
    (	253	)	,
    (	253	)	,
    (	253	)	,
    (	253	)	,
    (	253	)	,
    (	253	)	,
    (	253	)	,
    (	253	)	,
    (	252	)	,
    (	252	)	,
    (	252	)	,
    (	252	)	,
    (	252	)	,
    (	252	)	,
    (	252	)	,
    (	251	)	,
    (	251	)	,
    (	251	)	,
    (	251	)	,
    (	251	)	,
    (	251	)	,
    (	251	)	,
    (	250	)	,
    (	250	)	,
    (	250	)	,
    (	250	)	,
    (	250	)	,
    (	250	)	,
    (	250	)	,
    (	249	)	,
    (	249	)	,
    (	249	)	,
    (	249	)	,
    (	249	)	,
    (	249	)	,
    (	249	)	,
    (	249	)	,
    (	248	)	,
    (	248	)	,
    (	248	)	,
    (	248	)	,
    (	248	)	,
    (	248	)	,
    (	248	)	,
    (	247	)	,
    (	247	)	,
    (	247	)	,
    (	247	)	,
    (	247	)	,
    (	247	)	,
    (	247	)	,
    (	246	)	,
    (	246	)	,
    (	246	)	,
    (	246	)	,
    (	246	)	,
    (	246	)	,
    (	246	)	,
    (	245	)	,
    (	245	)	,
    (	245	)	,
    (	245	)	,
    (	245	)	,
    (	245	)	,
    (	245	)	,
    (	245	)	,
    (	244	)	,
    (	244	)	,
    (	244	)	,
    (	244	)	,
    (	244	)	,
    (	244	)	,
    (	244	)	,
    (	243	)	,
    (	243	)	,
    (	243	)	,
    (	243	)	,
    (	243	)	,
    (	243	)	,
    (	243	)	,
    (	242	)	,
    (	242	)	,
    (	242	)	,
    (	242	)	,
    (	242	)	,
    (	242	)	,
    (	242	)	,
    (	241	)	,
    (	241	)	,
    (	241	)	,
    (	241	)	,
    (	241	)	,
    (	241	)	,
    (	241	)	,
    (	241	)	,
    (	240	)	,
    (	240	)	,
    (	240	)	,
    (	240	)	,
    (	240	)	,
    (	240	)	,
    (	240	)	,
    (	239	)	,
    (	239	)	,
    (	239	)	,
    (	239	)	,
    (	239	)	,
    (	239	)	,
    (	239	)	,
    (	238	)	,
    (	238	)	,
    (	238	)	,
    (	238	)	,
    (	238	)	,
    (	238	)	,
    (	238	)	,
    (	237	)	,
    (	237	)	,
    (	237	)	,
    (	237	)	,
    (	237	)	,
    (	237	)	,
    (	237	)	,
    (	237	)	,
    (	236	)	,
    (	236	)	,
    (	236	)	,
    (	236	)	,
    (	236	)	,
    (	236	)	,
    (	236	)	,
    (	235	)	,
    (	235	)	,
    (	235	)	,
    (	235	)	,
    (	235	)	,
    (	235	)	,
    (	235	)	,
    (	234	)	,
    (	234	)	,
    (	234	)	,
    (	234	)	,
    (	234	)	,
    (	234	)	,
    (	234	)	,
    (	233	)	,
    (	233	)	,
    (	233	)	,
    (	233	)	,
    (	233	)	,
    (	233	)	,
    (	233	)	,
    (	233	)	,
    (	232	)	,
    (	232	)	,
    (	232	)	,
    (	232	)	,
    (	232	)	,
    (	232	)	,
    (	232	)	,
    (	231	)	,
    (	231	)	,
    (	231	)	,
    (	231	)	,
    (	231	)	,
    (	231	)	,
    (	231	)	,
    (	230	)	,
    (	230	)	,
    (	230	)	,
    (	230	)	,
    (	230	)	,
    (	230	)	,
    (	230	)	,
    (	229	)	,
    (	229	)	,
    (	229	)	,
    (	229	)	,
    (	229	)	,
    (	229	)	,
    (	229	)	,
    (	229	)	,
    (	228	)	,
    (	228	)	,
    (	228	)	,
    (	228	)	,
    (	228	)	,
    (	228	)	,
    (	228	)	,
    (	227	)	,
    (	227	)	,
    (	227	)	,
    (	227	)	,
    (	227	)	,
    (	227	)	,
    (	227	)	,
    (	226	)	,
    (	226	)	,
    (	226	)	,
    (	226	)	,
    (	226	)	,
    (	226	)	,
    (	226	)	,
    (	225	)	,
    (	225	)	,
    (	225	)	,
    (	225	)	,
    (	225	)	,
    (	225	)	,
    (	225	)	,
    (	225	)	,
    (	224	)	,
    (	224	)	,
    (	224	)	,
    (	224	)	,
    (	224	)	,
    (	224	)	,
    (	224	)	,
    (	223	)	,
    (	223	)	,
    (	223	)	,
    (	223	)	,
    (	223	)	,
    (	223	)	,
    (	223	)	,
    (	222	)	,
    (	222	)	,
    (	222	)	,
    (	222	)	,
    (	222	)	,
    (	222	)	,
    (	222	)	,
    (	221	)	,
    (	221	)	,
    (	221	)	,
    (	221	)	,
    (	221	)	,
    (	221	)	,
    (	221	)	,
    (	220	)	,
    (	220	)	,
    (	220	)	,
    (	220	)	,
    (	220	)	,
    (	220	)	,
    (	220	)	,
    (	220	)	,
    (	219	)	,
    (	219	)	,
    (	219	)	,
    (	219	)	,
    (	219	)	,
    (	219	)	,
    (	219	)	,
    (	218	)	,
    (	218	)	,
    (	218	)	,
    (	218	)	,
    (	218	)	,
    (	218	)	,
    (	218	)	,
    (	217	)	,
    (	217	)	,
    (	217	)	,
    (	217	)	,
    (	217	)	,
    (	217	)	,
    (	217	)	,
    (	216	)	,
    (	216	)	,
    (	216	)	,
    (	216	)	,
    (	216	)	,
    (	216	)	,
    (	216	)	,
    (	216	)	,
    (	215	)	,
    (	215	)	,
    (	215	)	,
    (	215	)	,
    (	215	)	,
    (	215	)	,
    (	215	)	,
    (	214	)	,
    (	214	)	,
    (	214	)	,
    (	214	)	,
    (	214	)	,
    (	214	)	,
    (	214	)	,
    (	213	)	,
    (	213	)	,
    (	213	)	,
    (	213	)	,
    (	213	)	,
    (	213	)	,
    (	213	)	,
    (	212	)	,
    (	212	)	,
    (	212	)	,
    (	212	)	,
    (	212	)	,
    (	212	)	,
    (	212	)	,
    (	212	)	,
    (	211	)	,
    (	211	)	,
    (	211	)	,
    (	211	)	,
    (	211	)	,
    (	211	)	,
    (	211	)	,
    (	210	)	,
    (	210	)	,
    (	210	)	,
    (	210	)	,
    (	210	)	,
    (	210	)	,
    (	210	)	,
    (	209	)	,
    (	209	)	,
    (	209	)	,
    (	209	)	,
    (	209	)	,
    (	209	)	,
    (	209	)	,
    (	208	)	,
    (	208	)	,
    (	208	)	,
    (	208	)	,
    (	208	)	,
    (	208	)	,
    (	208	)	,
    (	208	)	,
    (	207	)	,
    (	207	)	,
    (	207	)	,
    (	207	)	,
    (	207	)	,
    (	207	)	,
    (	207	)	,
    (	206	)	,
    (	206	)	,
    (	206	)	,
    (	206	)	,
    (	206	)	,
    (	206	)	,
    (	206	)	,
    (	205	)	,
    (	205	)	,
    (	205	)	,
    (	205	)	,
    (	205	)	,
    (	205	)	,
    (	205	)	,
    (	204	)	,
    (	204	)	,
    (	204	)	,
    (	204	)	,
    (	204	)	,
    (	204	)	,
    (	204	)	,
    (	204	)	,
    (	203	)	,
    (	203	)	,
    (	203	)	,
    (	203	)	,
    (	203	)	,
    (	203	)	,
    (	203	)	,
    (	202	)	,
    (	202	)	,
    (	202	)	,
    (	202	)	,
    (	202	)	,
    (	202	)	,
    (	202	)	,
    (	201	)	,
    (	201	)	,
    (	201	)	,
    (	201	)	,
    (	201	)	,
    (	201	)	,
    (	201	)	,
    (	200	)	,
    (	200	)	,
    (	200	)	,
    (	200	)	,
    (	200	)	,
    (	200	)	,
    (	200	)	,
    (	200	)	,
    (	199	)	,
    (	199	)	,
    (	199	)	,
    (	199	)	,
    (	199	)	,
    (	199	)	,
    (	199	)	,
    (	198	)	,
    (	198	)	,
    (	198	)	,
    (	198	)	,
    (	198	)	,
    (	198	)	,
    (	198	)	,
    (	197	)	,
    (	197	)	,
    (	197	)	,
    (	197	)	,
    (	197	)	,
    (	197	)	,
    (	197	)	,
    (	196	)	,
    (	196	)	,
    (	196	)	,
    (	196	)	,
    (	196	)	,
    (	196	)	,
    (	196	)	,
    (	196	)	,
    (	195	)	,
    (	195	)	,
    (	195	)	,
    (	195	)	,
    (	195	)	,
    (	195	)	,
    (	195	)	,
    (	194	)	,
    (	194	)	,
    (	194	)	,
    (	194	)	,
    (	194	)	,
    (	194	)	,
    (	194	)	,
    (	193	)	,
    (	193	)	,
    (	193	)	,
    (	193	)	,
    (	193	)	,
    (	193	)	,
    (	193	)	,
    (	192	)	,
    (	192	)	,
    (	192	)	,
    (	192	)	,
    (	192	)	,
    (	192	)	,
    (	192	)	,
    (	192	)	,
    (	191	)	,
    (	191	)	,
    (	191	)	,
    (	191	)	,
    (	191	)	,
    (	191	)	,
    (	191	)	,
    (	190	)	,
    (	190	)	,
    (	190	)	,
    (	190	)	,
    (	190	)	,
    (	190	)	,
    (	190	)	,
    (	189	)	,
    (	189	)	,
    (	189	)	,
    (	189	)	,
    (	189	)	,
    (	189	)	,
    (	189	)	,
    (	188	)	,
    (	188	)	,
    (	188	)	,
    (	188	)	,
    (	188	)	,
    (	188	)	,
    (	188	)	,
    (	188	)	,
    (	187	)	,
    (	187	)	,
    (	187	)	,
    (	187	)	,
    (	187	)	,
    (	187	)	,
    (	187	)	,
    (	186	)	,
    (	186	)	,
    (	186	)	,
    (	186	)	,
    (	186	)	,
    (	186	)	,
    (	186	)	,
    (	185	)	,
    (	185	)	,
    (	185	)	,
    (	185	)	,
    (	185	)	,
    (	185	)	,
    (	185	)	,
    (	184	)	,
    (	184	)	,
    (	184	)	,
    (	184	)	,
    (	184	)	,
    (	184	)	,
    (	184	)	,
    (	183	)	,
    (	183	)	,
    (	183	)	,
    (	183	)	,
    (	183	)	,
    (	183	)	,
    (	183	)	,
    (	183	)	,
    (	182	)	,
    (	182	)	,
    (	182	)	,
    (	182	)	,
    (	182	)	,
    (	182	)	,
    (	182	)	,
    (	181	)	,
    (	181	)	,
    (	181	)	,
    (	181	)	,
    (	181	)	,
    (	181	)	,
    (	181	)	,
    (	180	)	,
    (	180	)	,
    (	180	)	,
    (	180	)	,
    (	180	)	,
    (	180	)	,
    (	180	)	,
    (	179	)	,
    (	179	)	,
    (	179	)	,
    (	179	)	,
    (	179	)	,
    (	179	)	,
    (	179	)	,
    (	179	)	,
    (	178	)	,
    (	178	)	,
    (	178	)	,
    (	178	)	,
    (	178	)	,
    (	178	)	,
    (	178	)	,
    (	177	)	,
    (	177	)	,
    (	177	)	,
    (	177	)	,
    (	177	)	,
    (	177	)	,
    (	177	)	,
    (	176	)	,
    (	176	)	,
    (	176	)	,
    (	176	)	,
    (	176	)	,
    (	176	)	,
    (	176	)	,
    (	175	)	,
    (	175	)	,
    (	175	)	,
    (	175	)	,
    (	175	)	,
    (	175	)	,
    (	175	)	,
    (	175	)	,
    (	174	)	,
    (	174	)	,
    (	174	)	,
    (	174	)	,
    (	174	)	,
    (	174	)	,
    (	174	)	,
    (	173	)	,
    (	173	)	,
    (	173	)	,
    (	173	)	,
    (	173	)	,
    (	173	)	,
    (	173	)	,
    (	172	)	,
    (	172	)	,
    (	172	)	,
    (	172	)	,
    (	172	)	,
    (	172	)	,
    (	172	)	,
    (	171	)	,
    (	171	)	,
    (	171	)	,
    (	171	)	,
    (	171	)	,
    (	171	)	,
    (	171	)	,
    (	171	)	,
    (	170	)	,
    (	170	)	,
    (	170	)	,
    (	170	)	,
    (	170	)	,
    (	170	)	,
    (	170	)	,
    (	169	)	,
    (	169	)	,
    (	169	)	,
    (	169	)	,
    (	169	)	,
    (	169	)	,
    (	169	)	,
    (	168	)	,
    (	168	)	,
    (	168	)	,
    (	168	)	,
    (	168	)	,
    (	168	)	,
    (	168	)	,
    (	167	)	,
    (	167	)	,
    (	167	)	,
    (	167	)	,
    (	167	)	,
    (	167	)	,
    (	167	)	,
    (	167	)	,
    (	166	)	,
    (	166	)	,
    (	166	)	,
    (	166	)	,
    (	166	)	,
    (	166	)	,
    (	166	)	,
    (	165	)	,
    (	165	)	,
    (	165	)	,
    (	165	)	,
    (	165	)	,
    (	165	)	,
    (	165	)	,
    (	164	)	,
    (	164	)	,
    (	164	)	,
    (	164	)	,
    (	164	)	,
    (	164	)	,
    (	164	)	,
    (	163	)	,
    (	163	)	,
    (	163	)	,
    (	163	)	,
    (	163	)	,
    (	163	)	,
    (	163	)	,
    (	163	)	,
    (	162	)	,
    (	162	)	,
    (	162	)	,
    (	162	)	,
    (	162	)	,
    (	162	)	,
    (	162	)	,
    (	161	)	,
    (	161	)	,
    (	161	)	,
    (	161	)	,
    (	161	)	,
    (	161	)	,
    (	161	)	,
    (	160	)	,
    (	160	)	,
    (	160	)	,
    (	160	)	,
    (	160	)	,
    (	160	)	,
    (	160	)	,
    (	159	)	,
    (	159	)	,
    (	159	)	,
    (	159	)	,
    (	159	)	,
    (	159	)	,
    (	159	)	,
    (	159	)	,
    (	158	)	,
    (	158	)	,
    (	158	)	,
    (	158	)	,
    (	158	)	,
    (	158	)	,
    (	158	)	,
    (	157	)	,
    (	157	)	,
    (	157	)	,
    (	157	)	,
    (	157	)	,
    (	157	)	,
    (	157	)	,
    (	156	)	,
    (	156	)	,
    (	156	)	,
    (	156	)	,
    (	156	)	,
    (	156	)	,
    (	156	)	,
    (	155	)	,
    (	155	)	,
    (	155	)	,
    (	155	)	,
    (	155	)	,
    (	155	)	,
    (	155	)	,
    (	155	)	,
    (	154	)	,
    (	154	)	,
    (	154	)	,
    (	154	)	,
    (	154	)	,
    (	154	)	,
    (	154	)	,
    (	153	)	,
    (	153	)	,
    (	153	)	,
    (	153	)	,
    (	153	)	,
    (	153	)	,
    (	153	)	,
    (	152	)	,
    (	152	)	,
    (	152	)	,
    (	152	)	,
    (	152	)	,
    (	152	)	,
    (	152	)	,
    (	151	)	,
    (	151	)	,
    (	151	)	,
    (	151	)	,
    (	151	)	,
    (	151	)	,
    (	151	)	,
    (	150	)	,
    (	150	)	,
    (	150	)	,
    (	150	)	,
    (	150	)	,
    (	150	)	,
    (	150	)	,
    (	150	)	,
    (	149	)	,
    (	149	)	,
    (	149	)	,
    (	149	)	,
    (	149	)	,
    (	149	)	,
    (	149	)	,
    (	148	)	,
    (	148	)	,
    (	148	)	,
    (	148	)	,
    (	148	)	,
    (	148	)	,
    (	148	)	,
    (	147	)	,
    (	147	)	,
    (	147	)	,
    (	147	)	,
    (	147	)	,
    (	147	)	,
    (	147	)	,
    (	146	)	,
    (	146	)	,
    (	146	)	,
    (	146	)	,
    (	146	)	,
    (	146	)	,
    (	146	)	,
    (	146	)	,
    (	145	)	,
    (	145	)	,
    (	145	)	,
    (	145	)	,
    (	145	)	,
    (	145	)	,
    (	145	)	,
    (	144	)	,
    (	144	)	,
    (	144	)	,
    (	144	)	,
    (	144	)	,
    (	144	)	,
    (	144	)	,
    (	143	)	,
    (	143	)	,
    (	143	)	,
    (	143	)	,
    (	143	)	,
    (	143	)	,
    (	143	)	,
    (	142	)	,
    (	142	)	,
    (	142	)	,
    (	142	)	,
    (	142	)	,
    (	142	)	,
    (	142	)	,
    (	142	)	,
    (	141	)	,
    (	141	)	,
    (	141	)	,
    (	141	)	,
    (	141	)	,
    (	141	)	,
    (	141	)	,
    (	140	)	,
    (	140	)	,
    (	140	)	,
    (	140	)	,
    (	140	)	,
    (	140	)	,
    (	140	)	,
    (	139	)	,
    (	139	)	,
    (	139	)	,
    (	139	)	,
    (	139	)	,
    (	139	)	,
    (	139	)	,
    (	138	)	,
    (	138	)	,
    (	138	)	,
    (	138	)	,
    (	138	)	,
    (	138	)	,
    (	138	)	,
    (	138	)	,
    (	137	)	,
    (	137	)	,
    (	137	)	,
    (	137	)	,
    (	137	)	,
    (	137	)	,
    (	137	)	,
    (	136	)	,
    (	136	)	,
    (	136	)	,
    (	136	)	,
    (	136	)	,
    (	136	)	,
    (	136	)	,
    (	135	)	,
    (	135	)	,
    (	135	)	,
    (	135	)	,
    (	135	)	,
    (	135	)	,
    (	135	)	,
    (	134	)	,
    (	134	)	,
    (	134	)	,
    (	134	)	,
    (	134	)	,
    (	134	)	,
    (	134	)	,
    (	134	)	,
    (	133	)	,
    (	133	)	,
    (	133	)	,
    (	133	)	,
    (	133	)	,
    (	133	)	,
    (	133	)	,
    (	132	)	,
    (	132	)	,
    (	132	)	,
    (	132	)	,
    (	132	)	,
    (	132	)	,
    (	132	)	,
    (	131	)	,
    (	131	)	,
    (	131	)	,
    (	131	)	,
    (	131	)	,
    (	131	)	,
    (	131	)	,
    (	130	)	,
    (	130	)	,
    (	130	)	,
    (	130	)	,
    (	130	)	,
    (	130	)	,
    (	130	)	,
    (	130	)	,
    (	129	)	,
    (	129	)	,
    (	129	)	,
    (	129	)	,
    (	129	)	,
    (	129	)	,
    (	129	)	,
    (	128	)	,
    (	128	)	,
    (	128	)	,
    (	128	)	,
    (	128	)	,
    (	128	)	,
    (	128	)	,
    (	127	)	,
    (	127	)	,
    (	127	)	,
    (	127	)	,
    (	127	)	,
    (	127	)	,
    (	127	)	,
    (	126	)	,
    (	126	)	,
    (	126	)	,
    (	126	)	,
    (	126	)	,
    (	126	)	,
    (	126	)	,
    (	126	)	,
    (	125	)	,
    (	125	)	,
    (	125	)	,
    (	125	)	,
    (	125	)	,
    (	125	)	,
    (	125	)	,
    (	124	)	,
    (	124	)	,
    (	124	)	,
    (	124	)	,
    (	124	)	,
    (	124	)	,
    (	124	)	,
    (	123	)	,
    (	123	)	,
    (	123	)	,
    (	123	)	,
    (	123	)	,
    (	123	)	,
    (	123	)	,
    (	122	)	,
    (	122	)	,
    (	122	)	,
    (	122	)	,
    (	122	)	,
    (	122	)	,
    (	122	)	,
    (	122	)	,
    (	121	)	,
    (	121	)	,
    (	121	)	,
    (	121	)	,
    (	121	)	,
    (	121	)	,
    (	121	)	,
    (	120	)	,
    (	120	)	,
    (	120	)	,
    (	120	)	,
    (	120	)	,
    (	120	)	,
    (	120	)	,
    (	119	)	,
    (	119	)	,
    (	119	)	,
    (	119	)	,
    (	119	)	,
    (	119	)	,
    (	119	)	,
    (	118	)	,
    (	118	)	,
    (	118	)	,
    (	118	)	,
    (	118	)	,
    (	118	)	,
    (	118	)	,
    (	117	)	,
    (	117	)	,
    (	117	)	,
    (	117	)	,
    (	117	)	,
    (	117	)	,
    (	117	)	,
    (	117	)	,
    (	116	)	,
    (	116	)	,
    (	116	)	,
    (	116	)	,
    (	116	)	,
    (	116	)	,
    (	116	)	,
    (	115	)	,
    (	115	)	,
    (	115	)	,
    (	115	)	,
    (	115	)	,
    (	115	)	,
    (	115	)	,
    (	114	)	,
    (	114	)	,
    (	114	)	,
    (	114	)	,
    (	114	)	,
    (	114	)	,
    (	114	)	,
    (	113	)	,
    (	113	)	,
    (	113	)	,
    (	113	)	,
    (	113	)	,
    (	113	)	,
    (	113	)	,
    (	113	)	,
    (	112	)	,
    (	112	)	,
    (	112	)	,
    (	112	)	,
    (	112	)	,
    (	112	)	,
    (	112	)	,
    (	111	)	,
    (	111	)	,
    (	111	)	,
    (	111	)	,
    (	111	)	,
    (	111	)	,
    (	111	)	,
    (	110	)	,
    (	110	)	,
    (	110	)	,
    (	110	)	,
    (	110	)	,
    (	110	)	,
    (	110	)	,
    (	109	)	,
    (	109	)	,
    (	109	)	,
    (	109	)	,
    (	109	)	,
    (	109	)	,
    (	109	)	,
    (	109	)	,
    (	108	)	,
    (	108	)	,
    (	108	)	,
    (	108	)	,
    (	108	)	,
    (	108	)	,
    (	108	)	,
    (	107	)	,
    (	107	)	,
    (	107	)	,
    (	107	)	,
    (	107	)	,
    (	107	)	,
    (	107	)	,
    (	106	)	,
    (	106	)	,
    (	106	)	,
    (	106	)	,
    (	106	)	,
    (	106	)	,
    (	106	)	,
    (	105	)	,
    (	105	)	,
    (	105	)	,
    (	105	)	,
    (	105	)	,
    (	105	)	,
    (	105	)	,
    (	105	)	,
    (	104	)	,
    (	104	)	,
    (	104	)	,
    (	104	)	,
    (	104	)	,
    (	104	)	,
    (	104	)	,
    (	103	)	,
    (	103	)	,
    (	103	)	,
    (	103	)	,
    (	103	)	,
    (	103	)	,
    (	103	)	,
    (	102	)	,
    (	102	)	,
    (	102	)	,
    (	102	)	,
    (	102	)	,
    (	102	)	,
    (	102	)	,
    (	101	)	,
    (	101	)	,
    (	101	)	,
    (	101	)	,
    (	101	)	,
    (	101	)	,
    (	101	)	,
    (	101	)	,
    (	100	)	,
    (	100	)	,
    (	100	)	,
    (	100	)	,
    (	100	)	,
    (	100	)	,
    (	100	)	,
    (	99	)	,
    (	99	)	,
    (	99	)	,
    (	99	)	,
    (	99	)	,
    (	99	)	,
    (	99	)	,
    (	98	)	,
    (	98	)	,
    (	98	)	,
    (	98	)	,
    (	98	)	,
    (	98	)	,
    (	98	)	,
    (	97	)	,
    (	97	)	,
    (	97	)	,
    (	97	)	,
    (	97	)	,
    (	97	)	,
    (	97	)	,
    (	97	)	,
    (	96	)	,
    (	96	)	,
    (	96	)	,
    (	96	)	,
    (	96	)	,
    (	96	)	,
    (	96	)	,
    (	95	)	,
    (	95	)	,
    (	95	)	,
    (	95	)	,
    (	95	)	,
    (	95	)	,
    (	95	)	,
    (	94	)	,
    (	94	)	,
    (	94	)	,
    (	94	)	,
    (	94	)	,
    (	94	)	,
    (	94	)	,
    (	93	)	,
    (	93	)	,
    (	93	)	,
    (	93	)	,
    (	93	)	,
    (	93	)	,
    (	93	)	,
    (	93	)	,
    (	92	)	,
    (	92	)	,
    (	92	)	,
    (	92	)	,
    (	92	)	,
    (	92	)	,
    (	92	)	,
    (	91	)	,
    (	91	)	,
    (	91	)	,
    (	91	)	,
    (	91	)	,
    (	91	)	,
    (	91	)	,
    (	90	)	,
    (	90	)	,
    (	90	)	,
    (	90	)	,
    (	90	)	,
    (	90	)	,
    (	90	)	,
    (	89	)	,
    (	89	)	,
    (	89	)	,
    (	89	)	,
    (	89	)	,
    (	89	)	,
    (	89	)	,
    (	89	)	,
    (	88	)	,
    (	88	)	,
    (	88	)	,
    (	88	)	,
    (	88	)	,
    (	88	)	,
    (	88	)	,
    (	87	)	,
    (	87	)	,
    (	87	)	,
    (	87	)	,
    (	87	)	,
    (	87	)	,
    (	87	)	,
    (	86	)	,
    (	86	)	,
    (	86	)	,
    (	86	)	,
    (	86	)	,
    (	86	)	,
    (	86	)	,
    (	85	)	,
    (	85	)	,
    (	85	)	,
    (	85	)	,
    (	85	)	,
    (	85	)	,
    (	85	)	,
    (	84	)	,
    (	84	)	,
    (	84	)	,
    (	84	)	,
    (	84	)	,
    (	84	)	,
    (	84	)	,
    (	84	)	,
    (	83	)	,
    (	83	)	,
    (	83	)	,
    (	83	)	,
    (	83	)	,
    (	83	)	,
    (	83	)	,
    (	82	)	,
    (	82	)	,
    (	82	)	,
    (	82	)	,
    (	82	)	,
    (	82	)	,
    (	82	)	,
    (	81	)	,
    (	81	)	,
    (	81	)	,
    (	81	)	,
    (	81	)	,
    (	81	)	,
    (	81	)	,
    (	80	)	,
    (	80	)	,
    (	80	)	,
    (	80	)	,
    (	80	)	,
    (	80	)	,
    (	80	)	,
    (	80	)	,
    (	79	)	,
    (	79	)	,
    (	79	)	,
    (	79	)	,
    (	79	)	,
    (	79	)	,
    (	79	)	,
    (	78	)	,
    (	78	)	,
    (	78	)	,
    (	78	)	,
    (	78	)	,
    (	78	)	,
    (	78	)	,
    (	77	)	,
    (	77	)	,
    (	77	)	,
    (	77	)	,
    (	77	)	,
    (	77	)	,
    (	77	)	,
    (	76	)	,
    (	76	)	,
    (	76	)	,
    (	76	)	,
    (	76	)	,
    (	76	)	,
    (	76	)	,
    (	76	)	,
    (	75	)	,
    (	75	)	,
    (	75	)	,
    (	75	)	,
    (	75	)	,
    (	75	)	,
    (	75	)	,
    (	74	)	,
    (	74	)	,
    (	74	)	,
    (	74	)	,
    (	74	)	,
    (	74	)	,
    (	74	)	,
    (	73	)	,
    (	73	)	,
    (	73	)	,
    (	73	)	,
    (	73	)	,
    (	73	)	,
    (	73	)	,
    (	72	)	,
    (	72	)	,
    (	72	)	,
    (	72	)	,
    (	72	)	,
    (	72	)	,
    (	72	)	,
    (	72	)	,
    (	71	)	,
    (	71	)	,
    (	71	)	,
    (	71	)	,
    (	71	)	,
    (	71	)	,
    (	71	)	,
    (	70	)	,
    (	70	)	,
    (	70	)	,
    (	70	)	,
    (	70	)	,
    (	70	)	,
    (	70	)	,
    (	69	)	,
    (	69	)	,
    (	69	)	,
    (	69	)	,
    (	69	)	,
    (	69	)	,
    (	69	)	,
    (	68	)	,
    (	68	)	,
    (	68	)	,
    (	68	)	,
    (	68	)	,
    (	68	)	,
    (	68	)	,
    (	68	)	,
    (	67	)	,
    (	67	)	,
    (	67	)	,
    (	67	)	,
    (	67	)	,
    (	67	)	,
    (	67	)	,
    (	66	)	,
    (	66	)	,
    (	66	)	,
    (	66	)	,
    (	66	)	,
    (	66	)	,
    (	66	)	,
    (	65	)	,
    (	65	)	,
    (	65	)	,
    (	65	)	,
    (	65	)	,
    (	65	)	,
    (	65	)	,
    (	64	)	,
    (	64	)	,
    (	64	)	,
    (	64	)	,
    (	64	)	,
    (	64	)	,
    (	64	)	,
    (	64	)	,
    (	63	)	,
    (	63	)	,
    (	63	)	,
    (	63	)	,
    (	63	)	,
    (	63	)	,
    (	63	)	,
    (	62	)	,
    (	62	)	,
    (	62	)	,
    (	62	)	,
    (	62	)	,
    (	62	)	,
    (	62	)	,
    (	61	)	,
    (	61	)	,
    (	61	)	,
    (	61	)	,
    (	61	)	,
    (	61	)	,
    (	61	)	,
    (	60	)	,
    (	60	)	,
    (	60	)	,
    (	60	)	,
    (	60	)	,
    (	60	)	,
    (	60	)	,
    (	60	)	,
    (	59	)	,
    (	59	)	,
    (	59	)	,
    (	59	)	,
    (	59	)	,
    (	59	)	,
    (	59	)	,
    (	58	)	,
    (	58	)	,
    (	58	)	,
    (	58	)	,
    (	58	)	,
    (	58	)	,
    (	58	)	,
    (	57	)	,
    (	57	)	,
    (	57	)	,
    (	57	)	,
    (	57	)	,
    (	57	)	,
    (	57	)	,
    (	56	)	,
    (	56	)	,
    (	56	)	,
    (	56	)	,
    (	56	)	,
    (	56	)	,
    (	56	)	,
    (	56	)	,
    (	55	)	,
    (	55	)	,
    (	55	)	,
    (	55	)	,
    (	55	)	,
    (	55	)	,
    (	55	)	,
    (	54	)	,
    (	54	)	,
    (	54	)	,
    (	54	)	,
    (	54	)	,
    (	54	)	,
    (	54	)	,
    (	53	)	,
    (	53	)	,
    (	53	)	,
    (	53	)	,
    (	53	)	,
    (	53	)	,
    (	53	)	,
    (	52	)	,
    (	52	)	,
    (	52	)	,
    (	52	)	,
    (	52	)	,
    (	52	)	,
    (	52	)	,
    (	52	)	,
    (	51	)	,
    (	51	)	,
    (	51	)	,
    (	51	)	,
    (	51	)	,
    (	51	)	,
    (	51	)	,
    (	50	)	,
    (	50	)	,
    (	50	)	,
    (	50	)	,
    (	50	)	,
    (	50	)	,
    (	50	)	,
    (	49	)	,
    (	49	)	,
    (	49	)	,
    (	49	)	,
    (	49	)	,
    (	49	)	,
    (	49	)	,
    (	48	)	,
    (	48	)	,
    (	48	)	,
    (	48	)	,
    (	48	)	,
    (	48	)	,
    (	48	)	,
    (	47	)	,
    (	47	)	,
    (	47	)	,
    (	47	)	,
    (	47	)	,
    (	47	)	,
    (	47	)	,
    (	47	)	,
    (	46	)	,
    (	46	)	,
    (	46	)	,
    (	46	)	,
    (	46	)	,
    (	46	)	,
    (	46	)	,
    (	45	)	,
    (	45	)	,
    (	45	)	,
    (	45	)	,
    (	45	)	,
    (	45	)	,
    (	45	)	,
    (	44	)	,
    (	44	)	,
    (	44	)	,
    (	44	)	,
    (	44	)	,
    (	44	)	,
    (	44	)	,
    (	43	)	,
    (	43	)	,
    (	43	)	,
    (	43	)	,
    (	43	)	,
    (	43	)	,
    (	43	)	,
    (	43	)	,
    (	42	)	,
    (	42	)	,
    (	42	)	,
    (	42	)	,
    (	42	)	,
    (	42	)	,
    (	42	)	,
    (	41	)	,
    (	41	)	,
    (	41	)	,
    (	41	)	,
    (	41	)	,
    (	41	)	,
    (	41	)	,
    (	40	)	,
    (	40	)	,
    (	40	)	,
    (	40	)	,
    (	40	)	,
    (	40	)	,
    (	40	)	,
    (	39	)	,
    (	39	)	,
    (	39	)	,
    (	39	)	,
    (	39	)	,
    (	39	)	,
    (	39	)	,
    (	39	)	,
    (	38	)	,
    (	38	)	,
    (	38	)	,
    (	38	)	,
    (	38	)	,
    (	38	)	,
    (	38	)	,
    (	37	)	,
    (	37	)	,
    (	37	)	,
    (	37	)	,
    (	37	)	,
    (	37	)	,
    (	37	)	,
    (	36	)	,
    (	36	)	,
    (	36	)	,
    (	36	)	,
    (	36	)	,
    (	36	)	,
    (	36	)	,
    (	35	)	,
    (	35	)	,
    (	35	)	,
    (	35	)	,
    (	35	)	,
    (	35	)	,
    (	35	)	,
    (	35	)	,
    (	34	)	,
    (	34	)	,
    (	34	)	,
    (	34	)	,
    (	34	)	,
    (	34	)	,
    (	34	)	,
    (	33	)	,
    (	33	)	,
    (	33	)	,
    (	33	)	,
    (	33	)	,
    (	33	)	,
    (	33	)	,
    (	32	)	,
    (	32	)	,
    (	32	)	,
    (	32	)	,
    (	32	)	,
    (	32	)	,
    (	32	)	,
    (	31	)	,
    (	31	)	,
    (	31	)	,
    (	31	)	,
    (	31	)	,
    (	31	)	,
    (	31	)	,
    (	31	)	,
    (	30	)	,
    (	30	)	,
    (	30	)	,
    (	30	)	,
    (	30	)	,
    (	30	)	,
    (	30	)	,
    (	29	)	,
    (	29	)	,
    (	29	)	,
    (	29	)	,
    (	29	)	,
    (	29	)	,
    (	29	)	,
    (	28	)	,
    (	28	)	,
    (	28	)	,
    (	28	)	,
    (	28	)	,
    (	28	)	,
    (	28	)	,
    (	27	)	,
    (	27	)	,
    (	27	)	,
    (	27	)	,
    (	27	)	,
    (	27	)	,
    (	27	)	,
    (	27	)	,
    (	26	)	,
    (	26	)	,
    (	26	)	,
    (	26	)	,
    (	26	)	,
    (	26	)	,
    (	26	)	,
    (	25	)	,
    (	25	)	,
    (	25	)	,
    (	25	)	,
    (	25	)	,
    (	25	)	,
    (	25	)	,
    (	24	)	,
    (	24	)	,
    (	24	)	,
    (	24	)	,
    (	24	)	,
    (	24	)	,
    (	24	)	,
    (	23	)	,
    (	23	)	,
    (	23	)	,
    (	23	)	,
    (	23	)	,
    (	23	)	,
    (	23	)	,
    (	23	)	,
    (	22	)	,
    (	22	)	,
    (	22	)	,
    (	22	)	,
    (	22	)	,
    (	22	)	,
    (	22	)	,
    (	21	)	,
    (	21	)	,
    (	21	)	,
    (	21	)	,
    (	21	)	,
    (	21	)	,
    (	21	)	,
    (	20	)	,
    (	20	)	,
    (	20	)	,
    (	20	)	,
    (	20	)	,
    (	20	)	,
    (	20	)	,
    (	19	)	,
    (	19	)	,
    (	19	)	,
    (	19	)	,
    (	19	)	,
    (	19	)	,
    (	19	)	,
    (	19	)	,
    (	18	)	,
    (	18	)	,
    (	18	)	,
    (	18	)	,
    (	18	)	,
    (	18	)	,
    (	18	)	,
    (	17	)	,
    (	17	)	,
    (	17	)	,
    (	17	)	,
    (	17	)	,
    (	17	)	,
    (	17	)	,
    (	16	)	,
    (	16	)	,
    (	16	)	,
    (	16	)	,
    (	16	)	,
    (	16	)	,
    (	16	)	,
    (	15	)	,
    (	15	)	,
    (	15	)	,
    (	15	)	,
    (	15	)	,
    (	15	)	,
    (	15	)	,
    (	14	)	,
    (	14	)	,
    (	14	)	,
    (	14	)	,
    (	14	)	,
    (	14	)	,
    (	14	)	,
    (	14	)	,
    (	13	)	,
    (	13	)	,
    (	13	)	,
    (	13	)	,
    (	13	)	,
    (	13	)	,
    (	13	)	,
    (	12	)	,
    (	12	)	,
    (	12	)	,
    (	12	)	,
    (	12	)	,
    (	12	)	,
    (	12	)	,
    (	11	)	,
    (	11	)	,
    (	11	)	,
    (	11	)	,
    (	11	)	,
    (	11	)	,
    (	11	)	,
    (	10	)	,
    (	10	)	,
    (	10	)	,
    (	10	)	,
    (	10	)	,
    (	10	)	,
    (	10	)	,
    (	10	)	,
    (	9	)	,
    (	9	)	,
    (	9	)	,
    (	9	)	,
    (	9	)	,
    (	9	)	,
    (	9	)	,
    (	8	)	,
    (	8	)	,
    (	8	)	,
    (	8	)	,
    (	8	)	,
    (	8	)	,
    (	8	)	,
    (	7	)	,
    (	7	)	,
    (	7	)	,
    (	7	)	,
    (	7	)	,
    (	7	)	,
    (	7	)	,
    (	6	)	,
    (	6	)	,
    (	6	)	,
    (	6	)	,
    (	6	)	,
    (	6	)	,
    (	6	)	,
    (	6	)	,
    (	5	)	,
    (	5	)	,
    (	5	)	,
    (	5	)	,
    (	5	)	,
    (	5	)	,
    (	5	)	,
    (	4	)	,
    (	4	)	,
    (	4	)	,
    (	4	)	,
    (	4	)	,
    (	4	)	,
    (	4	)	,
    (	3	)	,
    (	3	)	,
    (	3	)	,
    (	3	)	,
    (	3	)	,
    (	3	)	,
    (	3	)	,
    (	2	)	,
    (	2	)	,
    (	2	)	,
    (	2	)	,
    (	2	)	,
    (	2	)	,
    (	2	)	,
    (	2	)	,
    (	1	)	,
    (	1	)	,
    (	1	)	,
    (	1	)	,
    (	1	)	,
    (	1	)	,
    (	1	)	,
    (	0	)	,
    (	0	)	,
    (	0	)	,
    (	0	)	
);

end package LUT_ledr;
