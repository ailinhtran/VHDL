library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_flash is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant flash_lut : array_1d := (
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    20    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    21    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    22    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    23    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    24    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    25    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    26    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    27    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    28    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    29    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    30    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    31    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    32    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    33    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    34    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    35    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    36    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    37    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    38    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    39    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    40    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    41    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    42    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    43    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    44    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    45    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    46    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    47    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    48    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    49    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    50    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    51    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    52    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    53    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    54    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    55    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    56    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    57    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    58    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    59    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    60    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    61    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    62    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    63    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    64    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    65    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    66    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    67    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    68    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    69    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    70    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    71    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    72    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    73    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    74    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    75    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    76    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    77    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    78    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    79    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    80    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    ,
(    1    )    

);

end package LUT_flash;
