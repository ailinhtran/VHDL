library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4092	)	,
(	4085	)	,
(	4077	)	,
(	4069	)	,
(	4062	)	,
(	4054	)	,
(	4047	)	,
(	4039	)	,
(	4032	)	,
(	4024	)	,
(	4017	)	,
(	4009	)	,
(	4002	)	,
(	3994	)	,
(	3987	)	,
(	3979	)	,
(	3972	)	,
(	3964	)	,
(	3957	)	,
(	3950	)	,
(	3942	)	,
(	3935	)	,
(	3928	)	,
(	3920	)	,
(	3913	)	,
(	3906	)	,
(	3898	)	,
(	3891	)	,
(	3884	)	,
(	3877	)	,
(	3869	)	,
(	3862	)	,
(	3855	)	,
(	3848	)	,
(	3840	)	,
(	3833	)	,
(	3826	)	,
(	3819	)	,
(	3812	)	,
(	3805	)	,
(	3798	)	,
(	3791	)	,
(	3784	)	,
(	3776	)	,
(	3769	)	,
(	3762	)	,
(	3755	)	,
(	3748	)	,
(	3741	)	,
(	3734	)	,
(	3727	)	,
(	3720	)	,
(	3714	)	,
(	3707	)	,
(	3700	)	,
(	3693	)	,
(	3686	)	,
(	3679	)	,
(	3672	)	,
(	3665	)	,
(	3658	)	,
(	3652	)	,
(	3645	)	,
(	3638	)	,
(	3631	)	,
(	3625	)	,
(	3618	)	,
(	3611	)	,
(	3604	)	,
(	3598	)	,
(	3591	)	,
(	3584	)	,
(	3578	)	,
(	3571	)	,
(	3564	)	,
(	3558	)	,
(	3551	)	,
(	3544	)	,
(	3538	)	,
(	3531	)	,
(	3525	)	,
(	3518	)	,
(	3511	)	,
(	3505	)	,
(	3498	)	,
(	3492	)	,
(	3485	)	,
(	3479	)	,
(	3472	)	,
(	3466	)	,
(	3460	)	,
(	3453	)	,
(	3447	)	,
(	3440	)	,
(	3434	)	,
(	3427	)	,
(	3421	)	,
(	3415	)	,
(	3408	)	,
(	3402	)	,
(	3396	)	,
(	3389	)	,
(	3383	)	,
(	3377	)	,
(	3371	)	,
(	3364	)	,
(	3358	)	,
(	3352	)	,
(	3346	)	,
(	3339	)	,
(	3333	)	,
(	3327	)	,
(	3321	)	,
(	3315	)	,
(	3309	)	,
(	3302	)	,
(	3296	)	,
(	3290	)	,
(	3284	)	,
(	3278	)	,
(	3272	)	,
(	3266	)	,
(	3260	)	,
(	3254	)	,
(	3248	)	,
(	3242	)	,
(	3236	)	,
(	3230	)	,
(	3224	)	,
(	3218	)	,
(	3212	)	,
(	3206	)	,
(	3200	)	,
(	3194	)	,
(	3188	)	,
(	3182	)	,
(	3176	)	,
(	3170	)	,
(	3165	)	,
(	3159	)	,
(	3153	)	,
(	3147	)	,
(	3141	)	,
(	3135	)	,
(	3130	)	,
(	3124	)	,
(	3118	)	,
(	3112	)	,
(	3107	)	,
(	3101	)	,
(	3095	)	,
(	3089	)	,
(	3084	)	,
(	3078	)	,
(	3072	)	,
(	3067	)	,
(	3061	)	,
(	3055	)	,
(	3050	)	,
(	3044	)	,
(	3039	)	,
(	3033	)	,
(	3027	)	,
(	3022	)	,
(	3016	)	,
(	3011	)	,
(	3005	)	,
(	3000	)	,
(	2994	)	,
(	2989	)	,
(	2983	)	,
(	2978	)	,
(	2972	)	,
(	2967	)	,
(	2961	)	,
(	2956	)	,
(	2951	)	,
(	2945	)	,
(	2940	)	,
(	2934	)	,
(	2929	)	,
(	2924	)	,
(	2918	)	,
(	2913	)	,
(	2908	)	,
(	2902	)	,
(	2897	)	,
(	2892	)	,
(	2886	)	,
(	2881	)	,
(	2876	)	,
(	2871	)	,
(	2865	)	,
(	2860	)	,
(	2855	)	,
(	2850	)	,
(	2844	)	,
(	2839	)	,
(	2834	)	,
(	2829	)	,
(	2824	)	,
(	2819	)	,
(	2813	)	,
(	2808	)	,
(	2803	)	,
(	2798	)	,
(	2793	)	,
(	2788	)	,
(	2783	)	,
(	2778	)	,
(	2773	)	,
(	2768	)	,
(	2763	)	,
(	2758	)	,
(	2753	)	,
(	2748	)	,
(	2743	)	,
(	2738	)	,
(	2733	)	,
(	2728	)	,
(	2723	)	,
(	2718	)	,
(	2713	)	,
(	2708	)	,
(	2703	)	,
(	2698	)	,
(	2693	)	,
(	2688	)	,
(	2684	)	,
(	2679	)	,
(	2674	)	,
(	2669	)	,
(	2664	)	,
(	2659	)	,
(	2655	)	,
(	2650	)	,
(	2645	)	,
(	2640	)	,
(	2636	)	,
(	2631	)	,
(	2626	)	,
(	2621	)	,
(	2617	)	,
(	2612	)	,
(	2607	)	,
(	2603	)	,
(	2598	)	,
(	2593	)	,
(	2589	)	,
(	2584	)	,
(	2579	)	,
(	2575	)	,
(	2570	)	,
(	2565	)	,
(	2561	)	,
(	2556	)	,
(	2552	)	,
(	2547	)	,
(	2543	)	,
(	2538	)	,
(	2534	)	,
(	2529	)	,
(	2524	)	,
(	2520	)	,
(	2515	)	,
(	2511	)	,
(	2507	)	,
(	2502	)	,
(	2498	)	,
(	2493	)	,
(	2489	)	,
(	2484	)	,
(	2480	)	,
(	2475	)	,
(	2471	)	,
(	2467	)	,
(	2462	)	,
(	2458	)	,
(	2454	)	,
(	2449	)	,
(	2445	)	,
(	2441	)	,
(	2436	)	,
(	2432	)	,
(	2428	)	,
(	2423	)	,
(	2419	)	,
(	2415	)	,
(	2411	)	,
(	2406	)	,
(	2402	)	,
(	2398	)	,
(	2394	)	,
(	2389	)	,
(	2385	)	,
(	2381	)	,
(	2377	)	,
(	2373	)	,
(	2368	)	,
(	2364	)	,
(	2360	)	,
(	2356	)	,
(	2352	)	,
(	2348	)	,
(	2344	)	,
(	2340	)	,
(	2335	)	,
(	2331	)	,
(	2327	)	,
(	2323	)	,
(	2319	)	,
(	2315	)	,
(	2311	)	,
(	2307	)	,
(	2303	)	,
(	2299	)	,
(	2295	)	,
(	2291	)	,
(	2287	)	,
(	2283	)	,
(	2279	)	,
(	2275	)	,
(	2271	)	,
(	2267	)	,
(	2263	)	,
(	2259	)	,
(	2256	)	,
(	2252	)	,
(	2248	)	,
(	2244	)	,
(	2240	)	,
(	2236	)	,
(	2232	)	,
(	2228	)	,
(	2225	)	,
(	2221	)	,
(	2217	)	,
(	2213	)	,
(	2209	)	,
(	2205	)	,
(	2202	)	,
(	2198	)	,
(	2194	)	,
(	2190	)	,
(	2187	)	,
(	2183	)	,
(	2179	)	,
(	2175	)	,
(	2172	)	,
(	2168	)	,
(	2164	)	,
(	2161	)	,
(	2157	)	,
(	2153	)	,
(	2150	)	,
(	2146	)	,
(	2142	)	,
(	2139	)	,
(	2135	)	,
(	2131	)	,
(	2128	)	,
(	2124	)	,
(	2121	)	,
(	2117	)	,
(	2113	)	,
(	2110	)	,
(	2106	)	,
(	2103	)	,
(	2099	)	,
(	2096	)	,
(	2092	)	,
(	2089	)	,
(	2085	)	,
(	2082	)	,
(	2078	)	,
(	2075	)	,
(	2071	)	,
(	2068	)	,
(	2064	)	,
(	2061	)	,
(	2057	)	,
(	2054	)	,
(	2050	)	,
(	2047	)	,
(	2044	)	,
(	2040	)	,
(	2037	)	,
(	2033	)	,
(	2030	)	,
(	2027	)	,
(	2023	)	,
(	2020	)	,
(	2017	)	,
(	2013	)	,
(	2010	)	,
(	2007	)	,
(	2003	)	,
(	2000	)	,
(	1997	)	,
(	1993	)	,
(	1990	)	,
(	1987	)	,
(	1984	)	,
(	1980	)	,
(	1977	)	,
(	1974	)	,
(	1971	)	,
(	1967	)	,
(	1964	)	,
(	1961	)	,
(	1958	)	,
(	1955	)	,
(	1951	)	,
(	1948	)	,
(	1945	)	,
(	1942	)	,
(	1939	)	,
(	1935	)	,
(	1932	)	,
(	1929	)	,
(	1926	)	,
(	1923	)	,
(	1920	)	,
(	1917	)	,
(	1914	)	,
(	1911	)	,
(	1907	)	,
(	1904	)	,
(	1901	)	,
(	1898	)	,
(	1895	)	,
(	1892	)	,
(	1889	)	,
(	1886	)	,
(	1883	)	,
(	1880	)	,
(	1877	)	,
(	1874	)	,
(	1871	)	,
(	1868	)	,
(	1865	)	,
(	1862	)	,
(	1859	)	,
(	1856	)	,
(	1853	)	,
(	1850	)	,
(	1847	)	,
(	1844	)	,
(	1842	)	,
(	1839	)	,
(	1836	)	,
(	1833	)	,
(	1830	)	,
(	1827	)	,
(	1824	)	,
(	1821	)	,
(	1818	)	,
(	1816	)	,
(	1813	)	,
(	1810	)	,
(	1807	)	,
(	1804	)	,
(	1801	)	,
(	1799	)	,
(	1796	)	,
(	1793	)	,
(	1790	)	,
(	1788	)	,
(	1785	)	,
(	1782	)	,
(	1779	)	,
(	1776	)	,
(	1774	)	,
(	1771	)	,
(	1768	)	,
(	1766	)	,
(	1763	)	,
(	1760	)	,
(	1757	)	,
(	1755	)	,
(	1752	)	,
(	1749	)	,
(	1747	)	,
(	1744	)	,
(	1741	)	,
(	1739	)	,
(	1736	)	,
(	1733	)	,
(	1731	)	,
(	1728	)	,
(	1725	)	,
(	1723	)	,
(	1720	)	,
(	1718	)	,
(	1715	)	,
(	1712	)	,
(	1710	)	,
(	1707	)	,
(	1705	)	,
(	1702	)	,
(	1700	)	,
(	1697	)	,
(	1695	)	,
(	1692	)	,
(	1689	)	,
(	1687	)	,
(	1684	)	,
(	1682	)	,
(	1679	)	,
(	1677	)	,
(	1674	)	,
(	1672	)	,
(	1669	)	,
(	1667	)	,
(	1665	)	,
(	1662	)	,
(	1660	)	,
(	1657	)	,
(	1655	)	,
(	1652	)	,
(	1650	)	,
(	1648	)	,
(	1645	)	,
(	1643	)	,
(	1640	)	,
(	1638	)	,
(	1636	)	,
(	1633	)	,
(	1631	)	,
(	1628	)	,
(	1626	)	,
(	1624	)	,
(	1621	)	,
(	1619	)	,
(	1617	)	,
(	1614	)	,
(	1612	)	,
(	1610	)	,
(	1607	)	,
(	1605	)	,
(	1603	)	,
(	1601	)	,
(	1598	)	,
(	1596	)	,
(	1594	)	,
(	1591	)	,
(	1589	)	,
(	1587	)	,
(	1585	)	,
(	1582	)	,
(	1580	)	,
(	1578	)	,
(	1576	)	,
(	1573	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1565	)	,
(	1562	)	,
(	1560	)	,
(	1558	)	,
(	1556	)	,
(	1554	)	,
(	1552	)	,
(	1549	)	,
(	1547	)	,
(	1545	)	,
(	1543	)	,
(	1541	)	,
(	1539	)	,
(	1537	)	,
(	1535	)	,
(	1532	)	,
(	1530	)	,
(	1528	)	,
(	1526	)	,
(	1524	)	,
(	1522	)	,
(	1520	)	,
(	1518	)	,
(	1516	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1508	)	,
(	1506	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1494	)	,
(	1492	)	,
(	1490	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1482	)	,
(	1480	)	,
(	1478	)	,
(	1476	)	,
(	1474	)	,
(	1472	)	,
(	1470	)	,
(	1468	)	,
(	1466	)	,
(	1464	)	,
(	1462	)	,
(	1460	)	,
(	1459	)	,
(	1457	)	,
(	1455	)	,
(	1453	)	,
(	1451	)	,
(	1449	)	,
(	1447	)	,
(	1445	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1433	)	,
(	1431	)	,
(	1429	)	,
(	1427	)	,
(	1425	)	,
(	1423	)	,
(	1422	)	,
(	1420	)	,
(	1418	)	,
(	1416	)	,
(	1415	)	,
(	1413	)	,
(	1411	)	,
(	1409	)	,
(	1407	)	,
(	1406	)	,
(	1404	)	,
(	1402	)	,
(	1401	)	,
(	1399	)	,
(	1397	)	,
(	1395	)	,
(	1394	)	,
(	1392	)	,
(	1390	)	,
(	1389	)	,
(	1387	)	,
(	1385	)	,
(	1383	)	,
(	1382	)	,
(	1380	)	,
(	1378	)	,
(	1377	)	,
(	1375	)	,
(	1373	)	,
(	1372	)	,
(	1370	)	,
(	1369	)	,
(	1367	)	,
(	1365	)	,
(	1364	)	,
(	1362	)	,
(	1360	)	,
(	1359	)	,
(	1357	)	,
(	1356	)	,
(	1354	)	,
(	1352	)	,
(	1351	)	,
(	1349	)	,
(	1348	)	,
(	1346	)	,
(	1345	)	,
(	1343	)	,
(	1341	)	,
(	1340	)	,
(	1338	)	,
(	1337	)	,
(	1335	)	,
(	1334	)	,
(	1332	)	,
(	1331	)	,
(	1329	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1323	)	,
(	1322	)	,
(	1320	)	,
(	1319	)	,
(	1317	)	,
(	1316	)	,
(	1314	)	,
(	1313	)	,
(	1311	)	,
(	1310	)	,
(	1308	)	,
(	1307	)	,
(	1305	)	,
(	1304	)	,
(	1302	)	,
(	1301	)	,
(	1300	)	,
(	1298	)	,
(	1297	)	,
(	1295	)	,
(	1294	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1288	)	,
(	1287	)	,
(	1286	)	,
(	1284	)	,
(	1283	)	,
(	1281	)	,
(	1280	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1275	)	,
(	1273	)	,
(	1272	)	,
(	1271	)	,
(	1269	)	,
(	1268	)	,
(	1266	)	,
(	1265	)	,
(	1264	)	,
(	1263	)	,
(	1261	)	,
(	1260	)	,
(	1259	)	,
(	1257	)	,
(	1256	)	,
(	1255	)	,
(	1253	)	,
(	1252	)	,
(	1251	)	,
(	1250	)	,
(	1248	)	,
(	1247	)	,
(	1246	)	,
(	1244	)	,
(	1243	)	,
(	1242	)	,
(	1241	)	,
(	1239	)	,
(	1238	)	,
(	1237	)	,
(	1236	)	,
(	1235	)	,
(	1233	)	,
(	1232	)	,
(	1231	)	,
(	1230	)	,
(	1228	)	,
(	1227	)	,
(	1226	)	,
(	1225	)	,
(	1224	)	,
(	1222	)	,
(	1221	)	,
(	1220	)	,
(	1219	)	,
(	1218	)	,
(	1216	)	,
(	1215	)	,
(	1214	)	,
(	1213	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1208	)	,
(	1207	)	,
(	1206	)	,
(	1205	)	,
(	1204	)	,
(	1203	)	,
(	1202	)	,
(	1200	)	,
(	1199	)	,
(	1198	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1192	)	,
(	1190	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1186	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1182	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1177	)	,
(	1176	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1165	)	,
(	1164	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1056	)	,
(	1055	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1049	)	,
(	1048	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1044	)	,
(	1043	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1041	)	,
(	1040	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1038	)	,
(	1037	)	,
(	1037	)	,
(	1036	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1034	)	,
(	1033	)	,
(	1033	)	,
(	1032	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1030	)	,
(	1029	)	,
(	1029	)	,
(	1028	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1026	)	,
(	1025	)	,
(	1025	)	,
(	1024	)	,
(	1024	)	,
(	1023	)	,
(	1023	)	,
(	1022	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1020	)	,
(	1019	)	,
(	1019	)	,
(	1018	)	,
(	1018	)	,
(	1017	)	,
(	1017	)	,
(	1016	)	,
(	1016	)	,
(	1015	)	,
(	1015	)	,
(	1014	)	,
(	1014	)	,
(	1013	)	,
(	1013	)	,
(	1012	)	,
(	1012	)	,
(	1011	)	,
(	1011	)	,
(	1010	)	,
(	1010	)	,
(	1009	)	,
(	1009	)	,
(	1008	)	,
(	1008	)	,
(	1007	)	,
(	1007	)	,
(	1006	)	,
(	1006	)	,
(	1005	)	,
(	1005	)	,
(	1004	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1002	)	,
(	1001	)	,
(	1001	)	,
(	1000	)	,
(	1000	)	,
(	1000	)	,
(	999	)	,
(	999	)	,
(	998	)	,
(	998	)	,
(	997	)	,
(	997	)	,
(	996	)	,
(	996	)	,
(	995	)	,
(	995	)	,
(	994	)	,
(	994	)	,
(	994	)	,
(	993	)	,
(	993	)	,
(	992	)	,
(	992	)	,
(	991	)	,
(	991	)	,
(	990	)	,
(	990	)	,
(	990	)	,
(	989	)	,
(	989	)	,
(	988	)	,
(	988	)	,
(	987	)	,
(	987	)	,
(	987	)	,
(	986	)	,
(	986	)	,
(	985	)	,
(	985	)	,
(	984	)	,
(	984	)	,
(	984	)	,
(	983	)	,
(	983	)	,
(	982	)	,
(	982	)	,
(	981	)	,
(	981	)	,
(	981	)	,
(	980	)	,
(	980	)	,
(	979	)	,
(	979	)	,
(	979	)	,
(	978	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	976	)	,
(	975	)	,
(	975	)	,
(	975	)	,
(	974	)	,
(	974	)	,
(	973	)	,
(	973	)	,
(	973	)	,
(	972	)	,
(	972	)	,
(	971	)	,
(	971	)	,
(	971	)	,
(	970	)	,
(	970	)	,
(	970	)	,
(	969	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	966	)	,
(	965	)	,
(	965	)	,
(	965	)	,
(	964	)	,
(	964	)	,
(	964	)	,
(	963	)	,
(	963	)	,
(	962	)	,
(	962	)	,
(	962	)	,
(	961	)	,
(	961	)	,
(	961	)	,
(	960	)	,
(	960	)	,
(	960	)	,
(	959	)	,
(	959	)	,
(	958	)	,
(	958	)	,
(	958	)	,
(	957	)	,
(	957	)	,
(	957	)	,
(	956	)	,
(	956	)	,
(	956	)	,
(	955	)	,
(	955	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	953	)	,
(	953	)	,
(	952	)	,
(	952	)	,
(	952	)	,
(	951	)	,
(	951	)	,
(	950	)	,
(	950	)	,
(	950	)	,
(	949	)	,
(	949	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	947	)	,
(	947	)	,
(	946	)	,
(	946	)	,
(	946	)	,
(	945	)	,
(	945	)	,
(	945	)	,
(	945	)	,
(	944	)	,
(	944	)	,
(	944	)	,
(	943	)	,
(	943	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	941	)	,
(	941	)	,
(	940	)	,
(	940	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	938	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	936	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	934	)	,
(	934	)	,
(	933	)	,
(	933	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	931	)	,
(	931	)	,
(	930	)	,
(	930	)	,
(	930	)	,
(	929	)	,
(	929	)	,
(	929	)	,
(	928	)	,
(	928	)	,
(	928	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	926	)	,
(	926	)	,
(	925	)	,
(	925	)	,
(	925	)	,
(	925	)	,
(	924	)	,
(	924	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	922	)	,
(	922	)	,
(	922	)	,
(	921	)	,
(	921	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	919	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	917	)	,
(	917	)	,
(	917	)	,
(	916	)	,
(	916	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	913	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	911	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	906	)	,
(	906	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	904	)	,
(	904	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	902	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	898	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	894	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	886	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	883	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	880	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	871	)	,
(	871	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	869	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	838	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	800	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	412	)	,
(	412	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	415	)	,
(	415	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	417	)	,
(	417	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	419	)	,
(	419	)	,
(	420	)	,
(	420	)	,
(	421	)	,
(	421	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	423	)	,
(	423	)	,
(	424	)	,
(	424	)	,
(	425	)	,
(	425	)	,
(	426	)	,
(	426	)	,
(	427	)	,
(	427	)	,
(	428	)	,
(	428	)	,
(	429	)	,
(	429	)	,
(	430	)	,
(	430	)	,
(	431	)	,
(	432	)	,
(	432	)	,
(	433	)	,
(	433	)	,
(	434	)	,
(	434	)	,
(	435	)	,
(	435	)	,
(	436	)	,
(	437	)	,
(	437	)	,
(	438	)	,
(	438	)	,
(	439	)	,
(	439	)	,
(	440	)	,
(	441	)	,
(	441	)	,
(	442	)	,
(	443	)	,
(	443	)	,
(	444	)	,
(	444	)	,
(	445	)	,
(	446	)	,
(	446	)	,
(	447	)	,
(	448	)	,
(	448	)	,
(	449	)	,
(	450	)	,
(	450	)	,
(	451	)	,
(	452	)	,
(	452	)	,
(	453	)	,
(	454	)	,
(	454	)	,
(	455	)	,
(	456	)	,
(	457	)	,
(	457	)	,
(	458	)	,
(	459	)	,
(	460	)	,
(	460	)	,
(	461	)	,
(	462	)	,
(	463	)	,
(	463	)	,
(	464	)	,
(	465	)	,
(	466	)	,
(	466	)	,
(	467	)	,
(	468	)	,
(	469	)	,
(	470	)	,
(	470	)	,
(	471	)	,
(	472	)	,
(	473	)	,
(	474	)	,
(	474	)	,
(	475	)	,
(	476	)	,
(	477	)	,
(	478	)	,
(	479	)	,
(	480	)	,
(	480	)	,
(	481	)	,
(	482	)	,
(	483	)	,
(	484	)	,
(	485	)	,
(	486	)	,
(	487	)	,
(	488	)	,
(	488	)	,
(	489	)	,
(	490	)	,
(	491	)	,
(	492	)	,
(	493	)	,
(	494	)	,
(	495	)	,
(	496	)	,
(	497	)	,
(	498	)	,
(	499	)	,
(	500	)	,
(	501	)	,
(	502	)	,
(	503	)	,
(	504	)	,
(	505	)	,
(	506	)	,
(	507	)	,
(	508	)	,
(	509	)	,
(	510	)	,
(	511	)	,
(	512	)	,
(	513	)	,
(	514	)	,
(	515	)	,
(	516	)	,
(	517	)	,
(	518	)	,
(	519	)	,
(	520	)	,
(	521	)	,
(	523	)	,
(	524	)	,
(	525	)	,
(	526	)	,
(	527	)	,
(	528	)	,
(	529	)	,
(	530	)	,
(	532	)	,
(	533	)	,
(	534	)	,
(	535	)	,
(	536	)	,
(	537	)	,
(	538	)	,
(	540	)	,
(	541	)	,
(	542	)	,
(	543	)	,
(	544	)	,
(	546	)	,
(	547	)	,
(	548	)	,
(	549	)	,
(	551	)	,
(	552	)	,
(	553	)	,
(	554	)	,
(	555	)	,
(	557	)	,
(	558	)	,
(	559	)	,
(	561	)	,
(	562	)	,
(	563	)	,
(	564	)	,
(	566	)	,
(	567	)	,
(	568	)	,
(	570	)	,
(	571	)	,
(	572	)	,
(	574	)	,
(	575	)	,
(	576	)	,
(	578	)	,
(	579	)	,
(	580	)	,
(	582	)	,
(	583	)	,
(	585	)	,
(	586	)	,
(	587	)	,
(	589	)	,
(	590	)	,
(	592	)	,
(	593	)	,
(	594	)	,
(	596	)	,
(	597	)	,
(	599	)	,
(	600	)	,
(	602	)	,
(	603	)	,
(	605	)	,
(	606	)	,
(	608	)	,
(	609	)	,
(	611	)	,
(	612	)	,
(	614	)	,
(	615	)	,
(	617	)	,
(	618	)	,
(	620	)	,
(	621	)	,
(	623	)	,
(	624	)	,
(	626	)	,
(	627	)	,
(	629	)	,
(	631	)	,
(	632	)	,
(	634	)	,
(	635	)	,
(	637	)	,
(	639	)	,
(	640	)	,
(	642	)	,
(	643	)	,
(	645	)	,
(	647	)	,
(	648	)	,
(	650	)	,
(	652	)	,
(	653	)	,
(	655	)	,
(	657	)	,
(	658	)	,
(	660	)	,
(	662	)	,
(	664	)	,
(	665	)	,
(	667	)	,
(	669	)	,
(	671	)	,
(	672	)	,
(	674	)	,
(	676	)	,
(	678	)	,
(	679	)	,
(	681	)	,
(	683	)	,
(	685	)	,
(	687	)	,
(	688	)	,
(	690	)	,
(	692	)	,
(	694	)	,
(	696	)	,
(	697	)	,
(	699	)	,
(	701	)	,
(	703	)	,
(	705	)	,
(	707	)	,
(	709	)	,
(	711	)	,
(	712	)	,
(	714	)	,
(	716	)	,
(	718	)	,
(	720	)	,
(	722	)	,
(	724	)	,
(	726	)	,
(	728	)	,
(	730	)	,
(	732	)	,
(	734	)	,
(	736	)	,
(	738	)	,
(	740	)	,
(	742	)	,
(	744	)	,
(	746	)	,
(	748	)	,
(	750	)	,
(	752	)	,
(	754	)	,
(	756	)	,
(	758	)	,
(	760	)	,
(	762	)	,
(	764	)	,
(	767	)	,
(	769	)	,
(	771	)	,
(	773	)	,
(	775	)	,
(	777	)	,
(	779	)	,
(	781	)	,
(	784	)	,
(	786	)	,
(	788	)	,
(	790	)	,
(	792	)	,
(	794	)	,
(	797	)	,
(	799	)	,
(	801	)	,
(	803	)	,
(	806	)	,
(	808	)	,
(	810	)	,
(	812	)	,
(	815	)	,
(	817	)	,
(	819	)	,
(	821	)	,
(	824	)	,
(	826	)	,
(	828	)	,
(	831	)	,
(	833	)	,
(	835	)	,
(	838	)	,
(	840	)	,
(	842	)	,
(	845	)	,
(	847	)	,
(	849	)	,
(	852	)	,
(	854	)	,
(	857	)	,
(	859	)	,
(	861	)	,
(	864	)	,
(	866	)	,
(	869	)	,
(	871	)	,
(	874	)	,
(	876	)	,
(	879	)	,
(	881	)	,
(	884	)	,
(	886	)	,
(	889	)	,
(	891	)	,
(	894	)	,
(	896	)	,
(	899	)	,
(	901	)	,
(	904	)	,
(	906	)	,
(	909	)	,
(	912	)	,
(	914	)	,
(	917	)	,
(	919	)	,
(	922	)	,
(	925	)	,
(	927	)	,
(	930	)	,
(	933	)	,
(	935	)	,
(	938	)	,
(	941	)	,
(	943	)	,
(	946	)	,
(	949	)	,
(	951	)	,
(	954	)	,
(	957	)	,
(	959	)	,
(	962	)	,
(	965	)	,
(	968	)	,
(	971	)	,
(	973	)	,
(	976	)	,
(	979	)	,
(	982	)	,
(	984	)	,
(	987	)	,
(	990	)	,
(	993	)	,
(	996	)	,
(	999	)	,
(	1002	)	,
(	1004	)	,
(	1007	)	,
(	1010	)	,
(	1013	)	,
(	1016	)	,
(	1019	)	,
(	1022	)	,
(	1025	)	,
(	1028	)	,
(	1031	)	,
(	1034	)	,
(	1037	)	,
(	1040	)	,
(	1043	)	,
(	1046	)	,
(	1049	)	,
(	1052	)	,
(	1055	)	,
(	1058	)	,
(	1061	)	,
(	1064	)	,
(	1067	)	,
(	1070	)	,
(	1073	)	,
(	1076	)	,
(	1079	)	,
(	1082	)	,
(	1085	)	,
(	1088	)	,
(	1092	)	,
(	1095	)	,
(	1098	)	,
(	1101	)	,
(	1104	)	,
(	1107	)	,
(	1111	)	,
(	1114	)	,
(	1117	)	,
(	1120	)	,
(	1123	)	,
(	1127	)	,
(	1130	)	,
(	1133	)	,
(	1136	)	,
(	1140	)	,
(	1143	)	,
(	1146	)	,
(	1150	)	,
(	1153	)	,
(	1156	)	,
(	1159	)	,
(	1163	)	,
(	1166	)	,
(	1170	)	,
(	1173	)	,
(	1176	)	,
(	1180	)	,
(	1183	)	,
(	1186	)	,
(	1190	)	,
(	1193	)	,
(	1197	)	,
(	1200	)	,
(	1204	)	,
(	1207	)	,
(	1211	)	,
(	1214	)	,
(	1217	)	,
(	1221	)	,
(	1225	)	,
(	1228	)	,
(	1232	)	,
(	1235	)	,
(	1239	)	,
(	1242	)	,
(	1246	)	,
(	1249	)	,
(	1253	)	,
(	1257	)	,
(	1260	)	,
(	1264	)	,
(	1267	)	,
(	1271	)	,
(	1275	)	,
(	1278	)	,
(	1282	)	,
(	1286	)	,
(	1289	)	,
(	1293	)	,
(	1297	)	,
(	1300	)	,
(	1304	)	,
(	1308	)	,
(	1312	)	,
(	1315	)	,
(	1319	)	,
(	1323	)	,
(	1327	)	,
(	1331	)	,
(	1334	)	,
(	1338	)	,
(	1342	)	,
(	1346	)	,
(	1350	)	,
(	1354	)	,
(	1357	)	,
(	1361	)	,
(	1365	)	,
(	1369	)	,
(	1373	)	,
(	1377	)	,
(	1381	)	,
(	1385	)	,
(	1389	)	,
(	1393	)	,
(	1397	)	,
(	1401	)	,
(	1405	)	,
(	1409	)	,
(	1413	)	,
(	1417	)	,
(	1421	)	,
(	1425	)	,
(	1429	)	,
(	1433	)	,
(	1437	)	,
(	1441	)	,
(	1445	)	,
(	1449	)	,
(	1453	)	,
(	1458	)	,
(	1462	)	,
(	1466	)	,
(	1470	)	,
(	1474	)	,
(	1478	)	,
(	1483	)	,
(	1487	)	,
(	1491	)	,
(	1495	)	,
(	1499	)	,
(	1504	)	,
(	1508	)	,
(	1512	)	,
(	1517	)	,
(	1521	)	,
(	1525	)	,
(	1529	)	,
(	1534	)	,
(	1538	)	,
(	1542	)	,
(	1547	)	,
(	1551	)	,
(	1556	)	,
(	1560	)	,
(	1564	)	,
(	1569	)	,
(	1573	)	,
(	1578	)	,
(	1582	)	,
(	1586	)	,
(	1591	)	,
(	1595	)	,
(	1600	)	,
(	1604	)	,
(	1609	)	,
(	1613	)	,
(	1618	)	,
(	1623	)	,
(	1627	)	,
(	1632	)	,
(	1636	)	,
(	1641	)	,
(	1645	)	,
(	1650	)	,
(	1655	)	,
(	1659	)	,
(	1664	)	,
(	1669	)	,
(	1673	)	,
(	1678	)	,
(	1683	)	,
(	1687	)	,
(	1692	)	,
(	1697	)	,
(	1702	)	,
(	1706	)	,
(	1711	)	,
(	1716	)	,
(	1721	)	,
(	1725	)	,
(	1730	)	,
(	1735	)	,
(	1740	)	,
(	1745	)	,
(	1750	)	,
(	1754	)	,
(	1759	)	,
(	1764	)	,
(	1769	)	,
(	1774	)	,
(	1779	)	,
(	1784	)	,
(	1789	)	,
(	1794	)	,
(	1799	)	,
(	1804	)	,
(	1809	)	,
(	1814	)	,
(	1819	)	,
(	1824	)	,
(	1829	)	,
(	1834	)	,
(	1839	)	,
(	1844	)	,
(	1849	)	,
(	1854	)	,
(	1859	)	,
(	1865	)	,
(	1870	)	,
(	1875	)	,
(	1880	)	,
(	1885	)	,
(	1890	)	,
(	1896	)	,
(	1901	)	,
(	1906	)	,
(	1911	)	,
(	1917	)	,
(	1922	)	,
(	1927	)	,
(	1932	)	,
(	1938	)	,
(	1943	)	,
(	1948	)	,
(	1954	)	,
(	1959	)	,
(	1964	)	,
(	1970	)	,
(	1975	)	,
(	1980	)	,
(	1986	)	,
(	1991	)	,
(	1997	)	,
(	2002	)	,
(	2008	)	,
(	2013	)	,
(	2019	)	,
(	2024	)	,
(	2030	)	,
(	2035	)	,
(	2041	)	,
(	2046	)	,
(	2052	)	,
(	2057	)	,
(	2063	)	,
(	2069	)	,
(	2074	)	,
(	2080	)	,
(	2085	)	,
(	2091	)	,
(	2097	)	,
(	2102	)	,
(	2108	)	,
(	2114	)	,
(	2119	)	,
(	2125	)	,
(	2131	)	,
(	2137	)	,
(	2142	)	,
(	2148	)	,
(	2154	)	,
(	2160	)	,
(	2166	)	,
(	2171	)	,
(	2177	)	,
(	2183	)	,
(	2189	)	,
(	2195	)	,
(	2201	)	,
(	2207	)	,
(	2213	)	,
(	2219	)	,
(	2225	)	,
(	2230	)	,
(	2236	)	,
(	2242	)	,
(	2248	)	,
(	2254	)	,
(	2260	)	,
(	2267	)	,
(	2273	)	,
(	2279	)	,
(	2285	)	,
(	2291	)	,
(	2297	)	,
(	2303	)	,
(	2309	)	,
(	2315	)	,
(	2321	)	,
(	2328	)	,
(	2334	)	,
(	2340	)	,
(	2346	)	,
(	2352	)	,
(	2359	)	,
(	2365	)	,
(	2371	)	,
(	2377	)	,
(	2384	)	,
(	2390	)	,
(	2396	)	,
(	2403	)	,
(	2409	)	,
(	2415	)	,
(	2422	)	,
(	2428	)	,
(	2435	)	,
(	2441	)	,
(	2447	)	,
(	2454	)	,
(	2460	)	,
(	2467	)	,
(	2473	)	,
(	2480	)	,
(	2486	)	,
(	2493	)	,
(	2499	)	,
(	2506	)	,
(	2513	)	,
(	2519	)	,
(	2526	)	,
(	2532	)	,
(	2539	)	,
(	2546	)	,
(	2552	)	,
(	2559	)	,
(	2566	)	,
(	2572	)	,
(	2579	)	,
(	2586	)	,
(	2592	)	,
(	2599	)	,
(	2606	)	,
(	2613	)	,
(	2620	)	,
(	2626	)	,
(	2633	)	,
(	2640	)	,
(	2647	)	,
(	2654	)	,
(	2661	)	,
(	2667	)	,
(	2674	)	,
(	2681	)	,
(	2688	)	,
(	2695	)	,
(	2702	)	,
(	2709	)	,
(	2716	)	,
(	2723	)	,
(	2730	)	,
(	2737	)	,
(	2744	)	,
(	2751	)	,
(	2758	)	,
(	2765	)	,
(	2773	)	,
(	2780	)	,
(	2787	)	,
(	2794	)	,
(	2801	)	,
(	2808	)	,
(	2816	)	,
(	2823	)	,
(	2830	)	,
(	2837	)	,
(	2845	)	,
(	2852	)	,
(	2859	)	,
(	2866	)	,
(	2874	)	,
(	2881	)	,
(	2888	)	,
(	2896	)	,
(	2903	)	,
(	2910	)	,
(	2918	)	,
(	2925	)	,
(	2933	)	,
(	2940	)	,
(	2948	)	,
(	2955	)	,
(	2963	)	,
(	2970	)	,
(	2978	)	,
(	2985	)	,
(	2993	)	,
(	3000	)	,
(	3008	)	,
(	3016	)	,
(	3023	)	,
(	3031	)	,
(	3038	)	,
(	3046	)	,
(	3054	)	,
(	3061	)	,
(	3069	)	,
(	3077	)	,
(	3085	)	,
(	3092	)	,
(	3100	)	,
(	3108	)	,
(	3116	)	,
(	3124	)	,
(	3131	)	,
(	3139	)	,
(	3147	)	,
(	3155	)	,
(	3163	)	,
(	3171	)	,
(	3179	)	,
(	3187	)	,
(	3195	)	,
(	3203	)	,
(	3211	)	,
(	3219	)	,
(	3227	)	,
(	3235	)	,
(	3243	)	,
(	3251	)	,
(	3259	)	,
(	3267	)	,
(	3275	)	,
(	3283	)	,
(	3291	)	,
(	3299	)	,
(	3308	)	,
(	3316	)	,
(	3324	)	,
(	3332	)	,
(	3340	)	,
(	3349	)	,
(	3357	)	,
(	3365	)	,
(	3374	)	,
(	3382	)	,
(	3390	)	,
(	3399	)	,
(	3407	)	,
(	3415	)	,
(	3424	)	,
(	3432	)	,
(	3441	)	,
(	3449	)	,
(	3457	)	,
(	3466	)	,
(	3474	)	,
(	3483	)	,
(	3492	)	,
(	3500	)	,
(	3509	)	,
(	3517	)	,
(	3526	)	,
(	3534	)	,
(	3543	)	,
(	3552	)	,
(	3560	)	,
(	3569	)	,
(	3578	)	,
(	3586	)	,
(	3595	)	,
(	3604	)	,
(	3613	)	,
(	3621	)	,
(	3630	)	,
(	3639	)	,
(	3648	)	,
(	3657	)	,
(	3666	)	,
(	3674	)	,
(	3683	)	,
(	3692	)	,
(	3701	)	,
(	3710	)	,
(	3719	)	,
(	3728	)	,
(	3737	)	,
(	3746	)	,
(	3755	)	,
(	3764	)	,
(	3773	)	,
(	3782	)	,
(	3791	)	,
(	3800	)	,
(	3810	)	,
(	3819	)	,
(	3828	)	,
(	3837	)	,
(	3846	)	,
(	3855	)	,
(	3865	)	,
(	3874	)	,
(	3883	)	,
(	3892	)	,
(	3902	)	,
(	3911	)	,
(	3920	)	,
(	3930	)	,
(	3939	)	,
(	3949	)	,
(	3958	)	,
(	3967	)	,
(	3977	)	,
(	3986	)	,
(	3996	)	,
(	4005	)	,
(	4015	)	,
(	4024	)	,
(	4034	)	,
(	4043	)	,
(	4053	)	,
(	4062	)	,
(	4072	)	,
(	4082	)	,
(	4091	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	    -- array index 4095 (voltage = "111111111111" or 4095 mV), distance output 3787 (37.87 cm)

);


end package LUT_pkg;
