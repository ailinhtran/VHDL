library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_flash is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant flash_lut : array_1d := (
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12500	)	,
(	12523	)	,
(	12547	)	,
(	12570	)	,
(	12593	)	,
(	12617	)	,
(	12640	)	,
(	12663	)	,
(	12687	)	,
(	12710	)	,
(	12733	)	,
(	12757	)	,
(	12780	)	,
(	12804	)	,
(	12827	)	,
(	12850	)	,
(	12874	)	,
(	12897	)	,
(	12920	)	,
(	12944	)	,
(	12967	)	,
(	12990	)	,
(	13014	)	,
(	13037	)	,
(	13060	)	,
(	13084	)	,
(	13107	)	,
(	13130	)	,
(	13154	)	,
(	13177	)	,
(	13200	)	,
(	13224	)	,
(	13247	)	,
(	13271	)	,
(	13294	)	,
(	13317	)	,
(	13341	)	,
(	13364	)	,
(	13387	)	,
(	13411	)	,
(	13434	)	,
(	13457	)	,
(	13481	)	,
(	13504	)	,
(	13527	)	,
(	13551	)	,
(	13574	)	,
(	13597	)	,
(	13621	)	,
(	13644	)	,
(	13667	)	,
(	13691	)	,
(	13714	)	,
(	13738	)	,
(	13761	)	,
(	13784	)	,
(	13808	)	,
(	13831	)	,
(	13854	)	,
(	13878	)	,
(	13901	)	,
(	13924	)	,
(	13948	)	,
(	13971	)	,
(	13994	)	,
(	14018	)	,
(	14041	)	,
(	14064	)	,
(	14088	)	,
(	14111	)	,
(	14134	)	,
(	14158	)	,
(	14181	)	,
(	14205	)	,
(	14228	)	,
(	14251	)	,
(	14275	)	,
(	14298	)	,
(	14321	)	,
(	14345	)	,
(	14368	)	,
(	14391	)	,
(	14415	)	,
(	14438	)	,
(	14461	)	,
(	14485	)	,
(	14508	)	,
(	14531	)	,
(	14555	)	,
(	14578	)	,
(	14601	)	,
(	14625	)	,
(	14648	)	,
(	14672	)	,
(	14695	)	,
(	14718	)	,
(	14742	)	,
(	14765	)	,
(	14788	)	,
(	14812	)	,
(	14835	)	,
(	14858	)	,
(	14882	)	,
(	14905	)	,
(	14928	)	,
(	14952	)	,
(	14975	)	,
(	14998	)	,
(	15022	)	,
(	15045	)	,
(	15068	)	,
(	15092	)	,
(	15115	)	,
(	15139	)	,
(	15162	)	,
(	15185	)	,
(	15209	)	,
(	15232	)	,
(	15255	)	,
(	15279	)	,
(	15302	)	,
(	15325	)	,
(	15349	)	,
(	15372	)	,
(	15395	)	,
(	15419	)	,
(	15442	)	,
(	15465	)	,
(	15489	)	,
(	15512	)	,
(	15535	)	,
(	15559	)	,
(	15582	)	,
(	15606	)	,
(	15629	)	,
(	15652	)	,
(	15676	)	,
(	15699	)	,
(	15722	)	,
(	15746	)	,
(	15769	)	,
(	15792	)	,
(	15816	)	,
(	15839	)	,
(	15862	)	,
(	15886	)	,
(	15909	)	,
(	15932	)	,
(	15956	)	,
(	15979	)	,
(	16002	)	,
(	16026	)	,
(	16049	)	,
(	16073	)	,
(	16096	)	,
(	16119	)	,
(	16143	)	,
(	16166	)	,
(	16189	)	,
(	16213	)	,
(	16236	)	,
(	16259	)	,
(	16283	)	,
(	16306	)	,
(	16329	)	,
(	16353	)	,
(	16376	)	,
(	16399	)	,
(	16423	)	,
(	16446	)	,
(	16469	)	,
(	16493	)	,
(	16516	)	,
(	16540	)	,
(	16563	)	,
(	16586	)	,
(	16610	)	,
(	16633	)	,
(	16656	)	,
(	16680	)	,
(	16703	)	,
(	16726	)	,
(	16750	)	,
(	16773	)	,
(	16796	)	,
(	16820	)	,
(	16843	)	,
(	16866	)	,
(	16890	)	,
(	16913	)	,
(	16936	)	,
(	16960	)	,
(	16983	)	,
(	17007	)	,
(	17030	)	,
(	17053	)	,
(	17077	)	,
(	17100	)	,
(	17123	)	,
(	17147	)	,
(	17170	)	,
(	17193	)	,
(	17217	)	,
(	17240	)	,
(	17263	)	,
(	17287	)	,
(	17310	)	,
(	17333	)	,
(	17357	)	,
(	17380	)	,
(	17403	)	,
(	17427	)	,
(	17450	)	,
(	17474	)	,
(	17497	)	,
(	17520	)	,
(	17544	)	,
(	17567	)	,
(	17590	)	,
(	17614	)	,
(	17637	)	,
(	17660	)	,
(	17684	)	,
(	17707	)	,
(	17730	)	,
(	17754	)	,
(	17777	)	,
(	17800	)	,
(	17824	)	,
(	17847	)	,
(	17870	)	,
(	17894	)	,
(	17917	)	,
(	17941	)	,
(	17964	)	,
(	17987	)	,
(	18011	)	,
(	18034	)	,
(	18057	)	,
(	18081	)	,
(	18104	)	,
(	18127	)	,
(	18151	)	,
(	18174	)	,
(	18197	)	,
(	18221	)	,
(	18244	)	,
(	18267	)	,
(	18291	)	,
(	18314	)	,
(	18337	)	,
(	18361	)	,
(	18384	)	,
(	18408	)	,
(	18431	)	,
(	18454	)	,
(	18478	)	,
(	18501	)	,
(	18524	)	,
(	18548	)	,
(	18571	)	,
(	18594	)	,
(	18618	)	,
(	18641	)	,
(	18664	)	,
(	18688	)	,
(	18711	)	,
(	18734	)	,
(	18758	)	,
(	18781	)	,
(	18804	)	,
(	18828	)	,
(	18851	)	,
(	18875	)	,
(	18898	)	,
(	18921	)	,
(	18945	)	,
(	18968	)	,
(	18991	)	,
(	19015	)	,
(	19038	)	,
(	19061	)	,
(	19085	)	,
(	19108	)	,
(	19131	)	,
(	19155	)	,
(	19178	)	,
(	19201	)	,
(	19225	)	,
(	19248	)	,
(	19271	)	,
(	19295	)	,
(	19318	)	,
(	19342	)	,
(	19365	)	,
(	19388	)	,
(	19412	)	,
(	19435	)	,
(	19458	)	,
(	19482	)	,
(	19505	)	,
(	19528	)	,
(	19552	)	,
(	19575	)	,
(	19598	)	,
(	19622	)	,
(	19645	)	,
(	19668	)	,
(	19692	)	,
(	19715	)	,
(	19738	)	,
(	19762	)	,
(	19785	)	,
(	19809	)	,
(	19832	)	,
(	19855	)	,
(	19879	)	,
(	19902	)	,
(	19925	)	,
(	19949	)	,
(	19972	)	,
(	19995	)	,
(	20019	)	,
(	20042	)	,
(	20065	)	,
(	20089	)	,
(	20112	)	,
(	20135	)	,
(	20159	)	,
(	20182	)	,
(	20205	)	,
(	20229	)	,
(	20252	)	,
(	20276	)	,
(	20299	)	,
(	20322	)	,
(	20346	)	,
(	20369	)	,
(	20392	)	,
(	20416	)	,
(	20439	)	,
(	20462	)	,
(	20486	)	,
(	20509	)	,
(	20532	)	,
(	20556	)	,
(	20579	)	,
(	20602	)	,
(	20626	)	,
(	20649	)	,
(	20672	)	,
(	20696	)	,
(	20719	)	,
(	20743	)	,
(	20766	)	,
(	20789	)	,
(	20813	)	,
(	20836	)	,
(	20859	)	,
(	20883	)	,
(	20906	)	,
(	20929	)	,
(	20953	)	,
(	20976	)	,
(	20999	)	,
(	21023	)	,
(	21046	)	,
(	21069	)	,
(	21093	)	,
(	21116	)	,
(	21139	)	,
(	21163	)	,
(	21186	)	,
(	21210	)	,
(	21233	)	,
(	21256	)	,
(	21280	)	,
(	21303	)	,
(	21326	)	,
(	21350	)	,
(	21373	)	,
(	21396	)	,
(	21420	)	,
(	21443	)	,
(	21466	)	,
(	21490	)	,
(	21513	)	,
(	21536	)	,
(	21560	)	,
(	21583	)	,
(	21606	)	,
(	21630	)	,
(	21653	)	,
(	21677	)	,
(	21700	)	,
(	21723	)	,
(	21747	)	,
(	21770	)	,
(	21793	)	,
(	21817	)	,
(	21840	)	,
(	21863	)	,
(	21887	)	,
(	21910	)	,
(	21933	)	,
(	21957	)	,
(	21980	)	,
(	22003	)	,
(	22027	)	,
(	22050	)	,
(	22073	)	,
(	22097	)	,
(	22120	)	,
(	22144	)	,
(	22167	)	,
(	22190	)	,
(	22214	)	,
(	22237	)	,
(	22260	)	,
(	22284	)	,
(	22307	)	,
(	22330	)	,
(	22354	)	,
(	22377	)	,
(	22400	)	,
(	22424	)	,
(	22447	)	,
(	22470	)	,
(	22494	)	,
(	22517	)	,
(	22540	)	,
(	22564	)	,
(	22587	)	,
(	22611	)	,
(	22634	)	,
(	22657	)	,
(	22681	)	,
(	22704	)	,
(	22727	)	,
(	22751	)	,
(	22774	)	,
(	22797	)	,
(	22821	)	,
(	22844	)	,
(	22867	)	,
(	22891	)	,
(	22914	)	,
(	22937	)	,
(	22961	)	,
(	22984	)	,
(	23007	)	,
(	23031	)	,
(	23054	)	,
(	23078	)	,
(	23101	)	,
(	23124	)	,
(	23148	)	,
(	23171	)	,
(	23194	)	,
(	23218	)	,
(	23241	)	,
(	23264	)	,
(	23288	)	,
(	23311	)	,
(	23334	)	,
(	23358	)	,
(	23381	)	,
(	23404	)	,
(	23428	)	,
(	23451	)	,
(	23474	)	,
(	23498	)	,
(	23521	)	,
(	23545	)	,
(	23568	)	,
(	23591	)	,
(	23615	)	,
(	23638	)	,
(	23661	)	,
(	23685	)	,
(	23708	)	,
(	23731	)	,
(	23755	)	,
(	23778	)	,
(	23801	)	,
(	23825	)	,
(	23848	)	,
(	23871	)	,
(	23895	)	,
(	23918	)	,
(	23941	)	,
(	23965	)	,
(	23988	)	,
(	24012	)	,
(	24035	)	,
(	24058	)	,
(	24082	)	,
(	24105	)	,
(	24128	)	,
(	24152	)	,
(	24175	)	,
(	24198	)	,
(	24222	)	,
(	24245	)	,
(	24268	)	,
(	24292	)	,
(	24315	)	,
(	24338	)	,
(	24362	)	,
(	24385	)	,
(	24408	)	,
(	24432	)	,
(	24455	)	,
(	24479	)	,
(	24502	)	,
(	24525	)	,
(	24549	)	,
(	24572	)	,
(	24595	)	,
(	24619	)	,
(	24642	)	,
(	24665	)	,
(	24689	)	,
(	24712	)	,
(	24735	)	,
(	24759	)	,
(	24782	)	,
(	24805	)	,
(	24829	)	,
(	24852	)	,
(	24875	)	,
(	24899	)	,
(	24922	)	,
(	24946	)	,
(	24969	)	,
(	24992	)	,
(	25016	)	,
(	25039	)	,
(	25062	)	,
(	25086	)	,
(	25109	)	,
(	25132	)	,
(	25156	)	,
(	25179	)	,
(	25202	)	,
(	25226	)	,
(	25249	)	,
(	25272	)	,
(	25296	)	,
(	25319	)	,
(	25342	)	,
(	25366	)	,
(	25389	)	,
(	25413	)	,
(	25436	)	,
(	25459	)	,
(	25483	)	,
(	25506	)	,
(	25529	)	,
(	25553	)	,
(	25576	)	,
(	25599	)	,
(	25623	)	,
(	25646	)	,
(	25669	)	,
(	25693	)	,
(	25716	)	,
(	25739	)	,
(	25763	)	,
(	25786	)	,
(	25809	)	,
(	25833	)	,
(	25856	)	,
(	25880	)	,
(	25903	)	,
(	25926	)	,
(	25950	)	,
(	25973	)	,
(	25996	)	,
(	26020	)	,
(	26043	)	,
(	26066	)	,
(	26090	)	,
(	26113	)	,
(	26136	)	,
(	26160	)	,
(	26183	)	,
(	26206	)	,
(	26230	)	,
(	26253	)	,
(	26276	)	,
(	26300	)	,
(	26323	)	,
(	26347	)	,
(	26370	)	,
(	26393	)	,
(	26417	)	,
(	26440	)	,
(	26463	)	,
(	26487	)	,
(	26510	)	,
(	26533	)	,
(	26557	)	,
(	26580	)	,
(	26603	)	,
(	26627	)	,
(	26650	)	,
(	26673	)	,
(	26697	)	,
(	26720	)	,
(	26743	)	,
(	26767	)	,
(	26790	)	,
(	26814	)	,
(	26837	)	,
(	26860	)	,
(	26884	)	,
(	26907	)	,
(	26930	)	,
(	26954	)	,
(	26977	)	,
(	27000	)	,
(	27024	)	,
(	27047	)	,
(	27070	)	,
(	27094	)	,
(	27117	)	,
(	27140	)	,
(	27164	)	,
(	27187	)	,
(	27210	)	,
(	27234	)	,
(	27257	)	,
(	27281	)	,
(	27304	)	,
(	27327	)	,
(	27351	)	,
(	27374	)	,
(	27397	)	,
(	27421	)	,
(	27444	)	,
(	27467	)	,
(	27491	)	,
(	27514	)	,
(	27537	)	,
(	27561	)	,
(	27584	)	,
(	27607	)	,
(	27631	)	,
(	27654	)	,
(	27677	)	,
(	27701	)	,
(	27724	)	,
(	27748	)	,
(	27771	)	,
(	27794	)	,
(	27818	)	,
(	27841	)	,
(	27864	)	,
(	27888	)	,
(	27911	)	,
(	27934	)	,
(	27958	)	,
(	27981	)	,
(	28004	)	,
(	28028	)	,
(	28051	)	,
(	28074	)	,
(	28098	)	,
(	28121	)	,
(	28144	)	,
(	28168	)	,
(	28191	)	,
(	28215	)	,
(	28238	)	,
(	28261	)	,
(	28285	)	,
(	28308	)	,
(	28331	)	,
(	28355	)	,
(	28378	)	,
(	28401	)	,
(	28425	)	,
(	28448	)	,
(	28471	)	,
(	28495	)	,
(	28518	)	,
(	28541	)	,
(	28565	)	,
(	28588	)	,
(	28611	)	,
(	28635	)	,
(	28658	)	,
(	28682	)	,
(	28705	)	,
(	28728	)	,
(	28752	)	,
(	28775	)	,
(	28798	)	,
(	28822	)	,
(	28845	)	,
(	28868	)	,
(	28892	)	,
(	28915	)	,
(	28938	)	,
(	28962	)	,
(	28985	)	,
(	29008	)	,
(	29032	)	,
(	29055	)	,
(	29078	)	,
(	29102	)	,
(	29125	)	,
(	29149	)	,
(	29172	)	,
(	29195	)	,
(	29219	)	,
(	29242	)	,
(	29265	)	,
(	29289	)	,
(	29312	)	,
(	29335	)	,
(	29359	)	,
(	29382	)	,
(	29405	)	,
(	29429	)	,
(	29452	)	,
(	29475	)	,
(	29499	)	,
(	29522	)	,
(	29545	)	,
(	29569	)	,
(	29592	)	,
(	29616	)	,
(	29639	)	,
(	29662	)	,
(	29686	)	,
(	29709	)	,
(	29732	)	,
(	29756	)	,
(	29779	)	,
(	29802	)	,
(	29826	)	,
(	29849	)	,
(	29872	)	,
(	29896	)	,
(	29919	)	,
(	29942	)	,
(	29966	)	,
(	29989	)	,
(	30012	)	,
(	30036	)	,
(	30059	)	,
(	30083	)	,
(	30106	)	,
(	30129	)	,
(	30153	)	,
(	30176	)	,
(	30199	)	,
(	30223	)	,
(	30246	)	,
(	30269	)	,
(	30293	)	,
(	30316	)	,
(	30339	)	,
(	30363	)	,
(	30386	)	,
(	30409	)	,
(	30433	)	,
(	30456	)	,
(	30479	)	,
(	30503	)	,
(	30526	)	,
(	30550	)	,
(	30573	)	,
(	30596	)	,
(	30620	)	,
(	30643	)	,
(	30666	)	,
(	30690	)	,
(	30713	)	,
(	30736	)	,
(	30760	)	,
(	30783	)	,
(	30806	)	,
(	30830	)	,
(	30853	)	,
(	30876	)	,
(	30900	)	,
(	30923	)	,
(	30946	)	,
(	30970	)	,
(	30993	)	,
(	31017	)	,
(	31040	)	,
(	31063	)	,
(	31087	)	,
(	31110	)	,
(	31133	)	,
(	31157	)	,
(	31180	)	,
(	31203	)	,
(	31227	)	,
(	31250	)	,
(	31273	)	,
(	31297	)	,
(	31320	)	,
(	31343	)	,
(	31367	)	,
(	31390	)	,
(	31413	)	,
(	31437	)	,
(	31460	)	,
(	31483	)	,
(	31507	)	,
(	31530	)	,
(	31554	)	,
(	31577	)	,
(	31600	)	,
(	31624	)	,
(	31647	)	,
(	31670	)	,
(	31694	)	,
(	31717	)	,
(	31740	)	,
(	31764	)	,
(	31787	)	,
(	31810	)	,
(	31834	)	,
(	31857	)	,
(	31880	)	,
(	31904	)	,
(	31927	)	,
(	31950	)	,
(	31974	)	,
(	31997	)	,
(	32021	)	,
(	32044	)	,
(	32067	)	,
(	32091	)	,
(	32114	)	,
(	32137	)	,
(	32161	)	,
(	32184	)	,
(	32207	)	,
(	32231	)	,
(	32254	)	,
(	32277	)	,
(	32301	)	,
(	32324	)	,
(	32347	)	,
(	32371	)	,
(	32394	)	,
(	32417	)	,
(	32441	)	,
(	32464	)	,
(	32488	)	,
(	32511	)	,
(	32534	)	,
(	32558	)	,
(	32581	)	,
(	32604	)	,
(	32628	)	,
(	32651	)	,
(	32674	)	,
(	32698	)	,
(	32721	)	,
(	32744	)	,
(	32768	)	,
(	32791	)	,
(	32814	)	,
(	32838	)	,
(	32861	)	,
(	32884	)	,
(	32908	)	,
(	32931	)	,
(	32955	)	,
(	32978	)	,
(	33001	)	,
(	33025	)	,
(	33048	)	,
(	33071	)	,
(	33095	)	,
(	33118	)	,
(	33141	)	,
(	33165	)	,
(	33188	)	,
(	33211	)	,
(	33235	)	,
(	33258	)	,
(	33281	)	,
(	33305	)	,
(	33328	)	,
(	33351	)	,
(	33375	)	,
(	33398	)	,
(	33422	)	,
(	33445	)	,
(	33468	)	,
(	33492	)	,
(	33515	)	,
(	33538	)	,
(	33562	)	,
(	33585	)	,
(	33608	)	,
(	33632	)	,
(	33655	)	,
(	33678	)	,
(	33702	)	,
(	33725	)	,
(	33748	)	,
(	33772	)	,
(	33795	)	,
(	33818	)	,
(	33842	)	,
(	33865	)	,
(	33889	)	,
(	33912	)	,
(	33935	)	,
(	33959	)	,
(	33982	)	,
(	34005	)	,
(	34029	)	,
(	34052	)	,
(	34075	)	,
(	34099	)	,
(	34122	)	,
(	34145	)	,
(	34169	)	,
(	34192	)	,
(	34215	)	,
(	34239	)	,
(	34262	)	,
(	34285	)	,
(	34309	)	,
(	34332	)	,
(	34356	)	,
(	34379	)	,
(	34402	)	,
(	34426	)	,
(	34449	)	,
(	34472	)	,
(	34496	)	,
(	34519	)	,
(	34542	)	,
(	34566	)	,
(	34589	)	,
(	34612	)	,
(	34636	)	,
(	34659	)	,
(	34682	)	,
(	34706	)	,
(	34729	)	,
(	34752	)	,
(	34776	)	,
(	34799	)	,
(	34823	)	,
(	34846	)	,
(	34869	)	,
(	34893	)	,
(	34916	)	,
(	34939	)	,
(	34963	)	,
(	34986	)	,
(	35009	)	,
(	35033	)	,
(	35056	)	,
(	35079	)	,
(	35103	)	,
(	35126	)	,
(	35149	)	,
(	35173	)	,
(	35196	)	,
(	35219	)	,
(	35243	)	,
(	35266	)	,
(	35290	)	,
(	35313	)	,
(	35336	)	,
(	35360	)	,
(	35383	)	,
(	35406	)	,
(	35430	)	,
(	35453	)	,
(	35476	)	,
(	35500	)	,
(	35523	)	,
(	35546	)	,
(	35570	)	,
(	35593	)	,
(	35616	)	,
(	35640	)	,
(	35663	)	,
(	35686	)	,
(	35710	)	,
(	35733	)	,
(	35757	)	,
(	35780	)	,
(	35803	)	,
(	35827	)	,
(	35850	)	,
(	35873	)	,
(	35897	)	,
(	35920	)	,
(	35943	)	,
(	35967	)	,
(	35990	)	,
(	36013	)	,
(	36037	)	,
(	36060	)	,
(	36083	)	,
(	36107	)	,
(	36130	)	,
(	36153	)	,
(	36177	)	,
(	36200	)	,
(	36224	)	,
(	36247	)	,
(	36270	)	,
(	36294	)	,
(	36317	)	,
(	36340	)	,
(	36364	)	,
(	36387	)	,
(	36410	)	,
(	36434	)	,
(	36457	)	,
(	36480	)	,
(	36504	)	,
(	36527	)	,
(	36550	)	,
(	36574	)	,
(	36597	)	,
(	36620	)	,
(	36644	)	,
(	36667	)	,
(	36691	)	,
(	36714	)	,
(	36737	)	,
(	36761	)	,
(	36784	)	,
(	36807	)	,
(	36831	)	,
(	36854	)	,
(	36877	)	,
(	36901	)	,
(	36924	)	,
(	36947	)	,
(	36971	)	,
(	36994	)	,
(	37017	)	,
(	37041	)	,
(	37064	)	,
(	37087	)	,
(	37111	)	,
(	37134	)	,
(	37158	)	,
(	37181	)	,
(	37204	)	,
(	37228	)	,
(	37251	)	,
(	37274	)	,
(	37298	)	,
(	37321	)	,
(	37344	)	,
(	37368	)	,
(	37391	)	,
(	37414	)	,
(	37438	)	,
(	37461	)	,
(	37484	)	,
(	37508	)	,
(	37531	)	,
(	37554	)	,
(	37578	)	,
(	37601	)	,
(	37625	)	,
(	37648	)	,
(	37671	)	,
(	37695	)	,
(	37718	)	,
(	37741	)	,
(	37765	)	,
(	37788	)	,
(	37811	)	,
(	37835	)	,
(	37858	)	,
(	37881	)	,
(	37905	)	,
(	37928	)	,
(	37951	)	,
(	37975	)	,
(	37998	)	,
(	38021	)	,
(	38045	)	,
(	38068	)	,
(	38092	)	,
(	38115	)	,
(	38138	)	,
(	38162	)	,
(	38185	)	,
(	38208	)	,
(	38232	)	,
(	38255	)	,
(	38278	)	,
(	38302	)	,
(	38325	)	,
(	38348	)	,
(	38372	)	,
(	38395	)	,
(	38418	)	,
(	38442	)	,
(	38465	)	,
(	38488	)	,
(	38512	)	,
(	38535	)	,
(	38559	)	,
(	38582	)	,
(	38605	)	,
(	38629	)	,
(	38652	)	,
(	38675	)	,
(	38699	)	,
(	38722	)	,
(	38745	)	,
(	38769	)	,
(	38792	)	,
(	38815	)	,
(	38839	)	,
(	38862	)	,
(	38885	)	,
(	38909	)	,
(	38932	)	,
(	38955	)	,
(	38979	)	,
(	39002	)	,
(	39026	)	,
(	39049	)	,
(	39072	)	,
(	39096	)	,
(	39119	)	,
(	39142	)	,
(	39166	)	,
(	39189	)	,
(	39212	)	,
(	39236	)	,
(	39259	)	,
(	39282	)	,
(	39306	)	,
(	39329	)	,
(	39352	)	,
(	39376	)	,
(	39399	)	,
(	39422	)	,
(	39446	)	,
(	39469	)	,
(	39493	)	,
(	39516	)	,
(	39539	)	,
(	39563	)	,
(	39586	)	,
(	39609	)	,
(	39633	)	,
(	39656	)	,
(	39679	)	,
(	39703	)	,
(	39726	)	,
(	39749	)	,
(	39773	)	,
(	39796	)	,
(	39819	)	,
(	39843	)	,
(	39866	)	,
(	39889	)	,
(	39913	)	,
(	39936	)	,
(	39960	)	,
(	39983	)	,
(	40006	)	,
(	40030	)	,
(	40053	)	,
(	40076	)	,
(	40100	)	,
(	40123	)	,
(	40146	)	,
(	40170	)	,
(	40193	)	,
(	40216	)	,
(	40240	)	,
(	40263	)	,
(	40286	)	,
(	40310	)	,
(	40333	)	,
(	40356	)	,
(	40380	)	,
(	40403	)	,
(	40427	)	,
(	40450	)	,
(	40473	)	,
(	40497	)	,
(	40520	)	,
(	40543	)	,
(	40567	)	,
(	40590	)	,
(	40613	)	,
(	40637	)	,
(	40660	)	,
(	40683	)	,
(	40707	)	,
(	40730	)	,
(	40753	)	,
(	40777	)	,
(	40800	)	,
(	40823	)	,
(	40847	)	,
(	40870	)	,
(	40894	)	,
(	40917	)	,
(	40940	)	,
(	40964	)	,
(	40987	)	,
(	41010	)	,
(	41034	)	,
(	41057	)	,
(	41080	)	,
(	41104	)	,
(	41127	)	,
(	41150	)	,
(	41174	)	,
(	41197	)	,
(	41220	)	,
(	41244	)	,
(	41267	)	,
(	41290	)	,
(	41314	)	,
(	41337	)	,
(	41361	)	,
(	41384	)	,
(	41407	)	,
(	41431	)	,
(	41454	)	,
(	41477	)	,
(	41501	)	,
(	41524	)	,
(	41547	)	,
(	41571	)	,
(	41594	)	,
(	41617	)	,
(	41641	)	,
(	41664	)	,
(	41687	)	,
(	41711	)	,
(	41734	)	,
(	41757	)	,
(	41781	)	,
(	41804	)	,
(	41828	)	,
(	41851	)	,
(	41874	)	,
(	41898	)	,
(	41921	)	,
(	41944	)	,
(	41968	)	,
(	41991	)	,
(	42014	)	,
(	42038	)	,
(	42061	)	,
(	42084	)	,
(	42108	)	,
(	42131	)	,
(	42154	)	,
(	42178	)	,
(	42201	)	,
(	42224	)	,
(	42248	)	,
(	42271	)	,
(	42295	)	,
(	42318	)	,
(	42341	)	,
(	42365	)	,
(	42388	)	,
(	42411	)	,
(	42435	)	,
(	42458	)	,
(	42481	)	,
(	42505	)	,
(	42528	)	,
(	42551	)	,
(	42575	)	,
(	42598	)	,
(	42621	)	,
(	42645	)	,
(	42668	)	,
(	42691	)	,
(	42715	)	,
(	42738	)	,
(	42762	)	,
(	42785	)	,
(	42808	)	,
(	42832	)	,
(	42855	)	,
(	42878	)	,
(	42902	)	,
(	42925	)	,
(	42948	)	,
(	42972	)	,
(	42995	)	,
(	43018	)	,
(	43042	)	,
(	43065	)	,
(	43088	)	,
(	43112	)	,
(	43135	)	,
(	43158	)	,
(	43182	)	,
(	43205	)	,
(	43229	)	,
(	43252	)	,
(	43275	)	,
(	43299	)	,
(	43322	)	,
(	43345	)	,
(	43369	)	,
(	43392	)	,
(	43415	)	,
(	43439	)	,
(	43462	)	,
(	43485	)	,
(	43509	)	,
(	43532	)	,
(	43555	)	,
(	43579	)	,
(	43602	)	,
(	43625	)	,
(	43649	)	,
(	43672	)	,
(	43696	)	,
(	43719	)	,
(	43742	)	,
(	43766	)	,
(	43789	)	,
(	43812	)	,
(	43836	)	,
(	43859	)	,
(	43882	)	,
(	43906	)	,
(	43929	)	,
(	43952	)	,
(	43976	)	,
(	43999	)	,
(	44022	)	,
(	44046	)	,
(	44069	)	,
(	44092	)	,
(	44116	)	,
(	44139	)	,
(	44163	)	,
(	44186	)	,
(	44209	)	,
(	44233	)	,
(	44256	)	,
(	44279	)	,
(	44303	)	,
(	44326	)	,
(	44349	)	,
(	44373	)	,
(	44396	)	,
(	44419	)	,
(	44443	)	,
(	44466	)	,
(	44489	)	,
(	44513	)	,
(	44536	)	,
(	44559	)	,
(	44583	)	,
(	44606	)	,
(	44630	)	,
(	44653	)	,
(	44676	)	,
(	44700	)	,
(	44723	)	,
(	44746	)	,
(	44770	)	,
(	44793	)	,
(	44816	)	,
(	44840	)	,
(	44863	)	,
(	44886	)	,
(	44910	)	,
(	44933	)	,
(	44956	)	,
(	44980	)	,
(	45003	)	,
(	45026	)	,
(	45050	)	,
(	45073	)	,
(	45097	)	,
(	45120	)	,
(	45143	)	,
(	45167	)	,
(	45190	)	,
(	45213	)	,
(	45237	)	,
(	45260	)	,
(	45283	)	,
(	45307	)	,
(	45330	)	,
(	45353	)	,
(	45377	)	,
(	45400	)	,
(	45423	)	,
(	45447	)	,
(	45470	)	,
(	45493	)	,
(	45517	)	,
(	45540	)	,
(	45564	)	,
(	45587	)	,
(	45610	)	,
(	45634	)	,
(	45657	)	,
(	45680	)	,
(	45704	)	,
(	45727	)	,
(	45750	)	,
(	45774	)	,
(	45797	)	,
(	45820	)	,
(	45844	)	,
(	45867	)	,
(	45890	)	,
(	45914	)	,
(	45937	)	,
(	45960	)	,
(	45984	)	,
(	46007	)	,
(	46031	)	,
(	46054	)	,
(	46077	)	,
(	46101	)	,
(	46124	)	,
(	46147	)	,
(	46171	)	,
(	46194	)	,
(	46217	)	,
(	46241	)	,
(	46264	)	,
(	46287	)	,
(	46311	)	,
(	46334	)	,
(	46357	)	,
(	46381	)	,
(	46404	)	,
(	46427	)	,
(	46451	)	,
(	46474	)	,
(	46498	)	,
(	46521	)	,
(	46544	)	,
(	46568	)	,
(	46591	)	,
(	46614	)	,
(	46638	)	,
(	46661	)	,
(	46684	)	,
(	46708	)	,
(	46731	)	,
(	46754	)	,
(	46778	)	,
(	46801	)	,
(	46824	)	,
(	46848	)	,
(	46871	)	,
(	46894	)	,
(	46918	)	,
(	46941	)	,
(	46965	)	,
(	46988	)	,
(	47011	)	,
(	47035	)	,
(	47058	)	,
(	47081	)	,
(	47105	)	,
(	47128	)	,
(	47151	)	,
(	47175	)	,
(	47198	)	,
(	47221	)	,
(	47245	)	,
(	47268	)	,
(	47291	)	,
(	47315	)	,
(	47338	)	,
(	47361	)	,
(	47385	)	,
(	47408	)	,
(	47432	)	,
(	47455	)	,
(	47478	)	,
(	47502	)	,
(	47525	)	,
(	47548	)	,
(	47572	)	,
(	47595	)	,
(	47618	)	,
(	47642	)	,
(	47665	)	,
(	47688	)	,
(	47712	)	,
(	47735	)	,
(	47758	)	,
(	47782	)	,
(	47805	)	,
(	47828	)	,
(	47852	)	,
(	47875	)	,
(	47899	)	,
(	47922	)	,
(	47945	)	,
(	47969	)	,
(	47992	)	,
(	48015	)	,
(	48039	)	,
(	48062	)	,
(	48085	)	,
(	48109	)	,
(	48132	)	,
(	48155	)	,
(	48179	)	,
(	48202	)	,
(	48225	)	,
(	48249	)	,
(	48272	)	,
(	48295	)	,
(	48319	)	,
(	48342	)	,
(	48366	)	,
(	48389	)	,
(	48412	)	,
(	48436	)	,
(	48459	)	,
(	48482	)	,
(	48506	)	,
(	48529	)	,
(	48552	)	,
(	48576	)	,
(	48599	)	,
(	48622	)	,
(	48646	)	,
(	48669	)	,
(	48692	)	,
(	48716	)	,
(	48739	)	,
(	48762	)	,
(	48786	)	,
(	48809	)	,
(	48833	)	,
(	48856	)	,
(	48879	)	,
(	48903	)	,
(	48926	)	,
(	48949	)	,
(	48973	)	,
(	48996	)	,
(	49019	)	,
(	49043	)	,
(	49066	)	,
(	49089	)	,
(	49113	)	,
(	49136	)	,
(	49159	)	,
(	49183	)	,
(	49206	)	,
(	49229	)	,
(	49253	)	,
(	49276	)	,
(	49300	)	,
(	49323	)	,
(	49346	)	,
(	49370	)	,
(	49393	)	,
(	49416	)	,
(	49440	)	,
(	49463	)	,
(	49486	)	,
(	49510	)	,
(	49533	)	,
(	49556	)	,
(	49580	)	,
(	49603	)	,
(	49626	)	,
(	49650	)	,
(	49673	)	,
(	49696	)	,
(	49720	)	,
(	49743	)	,
(	49767	)	,
(	49790	)	,
(	49813	)	,
(	49837	)	,
(	49860	)	,
(	49883	)	,
(	49907	)	,
(	49930	)	,
(	49953	)	,
(	49977	)	,
(	50000	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	

);

end package LUT_flash;
